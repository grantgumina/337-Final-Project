// $Id: $
// File name:   top.sv
// Created:     4/20/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: Top level file
