// $Id: $
// File name:   tb_usb_state_machine.sv
// Created:     4/16/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: Testbench for USB Protocol State Machine
