// $Id: $
// File name:   tb_datapath.sv
// Created:     4/16/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: Testbench for datapath block
