// $Id: $
// File name:   tb_usb_operation_controller.sv
// Created:     4/16/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: Testbench for usb operation controller
