
module bridge ( clk, n_rst, shift_en, data_in, data_out );
  input [7:0] data_in;
  output [511:0] data_out;
  input clk, n_rst, shift_en;
  wire   n523, n525, n527, n529, n531, n533, n535, n537, n539, n541, n543,
         n545, n547, n549, n551, n553, n555, n557, n559, n561, n563, n565,
         n567, n569, n571, n573, n575, n577, n579, n581, n583, n585, n587,
         n589, n591, n593, n595, n597, n599, n601, n603, n605, n607, n609,
         n611, n613, n615, n617, n619, n621, n623, n625, n627, n629, n631,
         n633, n635, n637, n639, n641, n643, n645, n647, n649, n651, n653,
         n655, n657, n659, n661, n663, n665, n667, n669, n671, n673, n675,
         n677, n679, n681, n683, n685, n687, n689, n691, n693, n695, n697,
         n699, n701, n703, n705, n707, n709, n711, n713, n715, n717, n719,
         n721, n723, n725, n727, n729, n731, n733, n735, n737, n739, n741,
         n743, n745, n747, n749, n751, n753, n755, n757, n759, n761, n763,
         n765, n767, n769, n771, n773, n775, n777, n779, n781, n783, n785,
         n787, n789, n791, n793, n795, n797, n799, n801, n803, n805, n807,
         n809, n811, n813, n815, n817, n819, n821, n823, n825, n827, n829,
         n831, n833, n835, n837, n839, n841, n843, n845, n847, n849, n851,
         n853, n855, n857, n859, n861, n863, n865, n867, n869, n871, n873,
         n875, n877, n879, n881, n883, n885, n887, n889, n891, n893, n895,
         n897, n899, n901, n903, n905, n907, n909, n911, n913, n915, n917,
         n919, n921, n923, n925, n927, n929, n931, n933, n935, n937, n939,
         n941, n943, n945, n947, n949, n951, n953, n955, n957, n959, n961,
         n963, n965, n967, n969, n971, n973, n975, n977, n979, n981, n983,
         n985, n987, n989, n991, n993, n995, n997, n999, n1001, n1003, n1005,
         n1007, n1009, n1011, n1013, n1015, n1017, n1019, n1021, n1023, n1025,
         n1027, n1029, n1031, n1033, n1035, n1037, n1039, n1041, n1043, n1045,
         n1047, n1049, n1051, n1053, n1055, n1057, n1059, n1061, n1063, n1065,
         n1067, n1069, n1071, n1073, n1075, n1077, n1079, n1081, n1083, n1085,
         n1087, n1089, n1091, n1093, n1095, n1097, n1099, n1101, n1103, n1105,
         n1107, n1109, n1111, n1113, n1115, n1117, n1119, n1121, n1123, n1125,
         n1127, n1129, n1131, n1133, n1135, n1137, n1139, n1141, n1143, n1145,
         n1147, n1149, n1151, n1153, n1155, n1157, n1159, n1161, n1163, n1165,
         n1167, n1169, n1171, n1173, n1175, n1177, n1179, n1181, n1183, n1185,
         n1187, n1189, n1191, n1193, n1195, n1197, n1199, n1201, n1203, n1205,
         n1207, n1209, n1211, n1213, n1215, n1217, n1219, n1221, n1223, n1225,
         n1227, n1229, n1231, n1233, n1235, n1237, n1239, n1241, n1243, n1245,
         n1247, n1249, n1251, n1253, n1255, n1257, n1259, n1261, n1263, n1265,
         n1267, n1269, n1271, n1273, n1275, n1277, n1279, n1281, n1283, n1285,
         n1287, n1289, n1291, n1293, n1295, n1297, n1299, n1301, n1303, n1305,
         n1307, n1309, n1311, n1313, n1315, n1317, n1319, n1321, n1323, n1325,
         n1327, n1329, n1331, n1333, n1335, n1337, n1339, n1341, n1343, n1345,
         n1347, n1349, n1351, n1353, n1355, n1357, n1359, n1361, n1363, n1365,
         n1367, n1369, n1371, n1373, n1375, n1377, n1379, n1381, n1383, n1385,
         n1387, n1389, n1391, n1393, n1395, n1397, n1399, n1401, n1403, n1405,
         n1407, n1409, n1411, n1413, n1415, n1417, n1419, n1421, n1423, n1425,
         n1427, n1429, n1431, n1433, n1435, n1437, n1439, n1441, n1443, n1445,
         n1447, n1449, n1451, n1453, n1455, n1457, n1459, n1461, n1463, n1465,
         n1467, n1469, n1471, n1473, n1475, n1477, n1479, n1481, n1483, n1485,
         n1487, n1489, n1491, n1493, n1495, n1497, n1499, n1501, n1503, n1505,
         n1507, n1509, n1511, n1513, n1515, n1517, n1519, n1521, n1523, n1525,
         n1527, n1529, n1531, n1533, n1535, n1537, n1539, n1541, n1543, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057;

  DFFSR \current_reg[7]  ( .D(n1545), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[7]) );
  DFFSR \current_reg[15]  ( .D(n1543), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[15]) );
  DFFSR \current_reg[23]  ( .D(n1541), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[23]) );
  DFFSR \current_reg[31]  ( .D(n1539), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[31]) );
  DFFSR \current_reg[39]  ( .D(n1537), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[39]) );
  DFFSR \current_reg[47]  ( .D(n1535), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[47]) );
  DFFSR \current_reg[55]  ( .D(n1533), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[55]) );
  DFFSR \current_reg[63]  ( .D(n1531), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[63]) );
  DFFSR \current_reg[71]  ( .D(n1529), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[71]) );
  DFFSR \current_reg[79]  ( .D(n1527), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[79]) );
  DFFSR \current_reg[87]  ( .D(n1525), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[87]) );
  DFFSR \current_reg[95]  ( .D(n1523), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[95]) );
  DFFSR \current_reg[103]  ( .D(n1521), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[103]) );
  DFFSR \current_reg[111]  ( .D(n1519), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[111]) );
  DFFSR \current_reg[119]  ( .D(n1517), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[119]) );
  DFFSR \current_reg[127]  ( .D(n1515), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[127]) );
  DFFSR \current_reg[135]  ( .D(n1513), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[135]) );
  DFFSR \current_reg[143]  ( .D(n1511), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[143]) );
  DFFSR \current_reg[151]  ( .D(n1509), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[151]) );
  DFFSR \current_reg[159]  ( .D(n1507), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[159]) );
  DFFSR \current_reg[167]  ( .D(n1505), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[167]) );
  DFFSR \current_reg[175]  ( .D(n1503), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[175]) );
  DFFSR \current_reg[183]  ( .D(n1501), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[183]) );
  DFFSR \current_reg[191]  ( .D(n1499), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[191]) );
  DFFSR \current_reg[199]  ( .D(n1497), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[199]) );
  DFFSR \current_reg[207]  ( .D(n1495), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[207]) );
  DFFSR \current_reg[215]  ( .D(n1493), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[215]) );
  DFFSR \current_reg[223]  ( .D(n1491), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[223]) );
  DFFSR \current_reg[231]  ( .D(n1489), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[231]) );
  DFFSR \current_reg[239]  ( .D(n1487), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[239]) );
  DFFSR \current_reg[247]  ( .D(n1485), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[247]) );
  DFFSR \current_reg[255]  ( .D(n1483), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[255]) );
  DFFSR \current_reg[263]  ( .D(n1481), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[263]) );
  DFFSR \current_reg[271]  ( .D(n1479), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[271]) );
  DFFSR \current_reg[279]  ( .D(n1477), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[279]) );
  DFFSR \current_reg[287]  ( .D(n1475), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[287]) );
  DFFSR \current_reg[295]  ( .D(n1473), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[295]) );
  DFFSR \current_reg[303]  ( .D(n1471), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[303]) );
  DFFSR \current_reg[311]  ( .D(n1469), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[311]) );
  DFFSR \current_reg[319]  ( .D(n1467), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[319]) );
  DFFSR \current_reg[327]  ( .D(n1465), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[327]) );
  DFFSR \current_reg[335]  ( .D(n1463), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[335]) );
  DFFSR \current_reg[343]  ( .D(n1461), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[343]) );
  DFFSR \current_reg[351]  ( .D(n1459), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[351]) );
  DFFSR \current_reg[359]  ( .D(n1457), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[359]) );
  DFFSR \current_reg[367]  ( .D(n1455), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[367]) );
  DFFSR \current_reg[375]  ( .D(n1453), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[375]) );
  DFFSR \current_reg[383]  ( .D(n1451), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[383]) );
  DFFSR \current_reg[391]  ( .D(n1449), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[391]) );
  DFFSR \current_reg[399]  ( .D(n1447), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[399]) );
  DFFSR \current_reg[407]  ( .D(n1445), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[407]) );
  DFFSR \current_reg[415]  ( .D(n1443), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[415]) );
  DFFSR \current_reg[423]  ( .D(n1441), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[423]) );
  DFFSR \current_reg[431]  ( .D(n1439), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[431]) );
  DFFSR \current_reg[439]  ( .D(n1437), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[439]) );
  DFFSR \current_reg[447]  ( .D(n1435), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[447]) );
  DFFSR \current_reg[455]  ( .D(n1433), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[455]) );
  DFFSR \current_reg[463]  ( .D(n1431), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[463]) );
  DFFSR \current_reg[471]  ( .D(n1429), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[471]) );
  DFFSR \current_reg[479]  ( .D(n1427), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[479]) );
  DFFSR \current_reg[487]  ( .D(n1425), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[487]) );
  DFFSR \current_reg[495]  ( .D(n1423), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[495]) );
  DFFSR \current_reg[503]  ( .D(n1421), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[503]) );
  DFFSR \current_reg[511]  ( .D(n1419), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[511]) );
  DFFSR \current_reg[6]  ( .D(n1417), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[6]) );
  DFFSR \current_reg[14]  ( .D(n1415), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[14]) );
  DFFSR \current_reg[22]  ( .D(n1413), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[22]) );
  DFFSR \current_reg[30]  ( .D(n1411), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[30]) );
  DFFSR \current_reg[38]  ( .D(n1409), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[38]) );
  DFFSR \current_reg[46]  ( .D(n1407), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[46]) );
  DFFSR \current_reg[54]  ( .D(n1405), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[54]) );
  DFFSR \current_reg[62]  ( .D(n1403), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[62]) );
  DFFSR \current_reg[70]  ( .D(n1401), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[70]) );
  DFFSR \current_reg[78]  ( .D(n1399), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[78]) );
  DFFSR \current_reg[86]  ( .D(n1397), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[86]) );
  DFFSR \current_reg[94]  ( .D(n1395), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[94]) );
  DFFSR \current_reg[102]  ( .D(n1393), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[102]) );
  DFFSR \current_reg[110]  ( .D(n1391), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[110]) );
  DFFSR \current_reg[118]  ( .D(n1389), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[118]) );
  DFFSR \current_reg[126]  ( .D(n1387), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[126]) );
  DFFSR \current_reg[134]  ( .D(n1385), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[134]) );
  DFFSR \current_reg[142]  ( .D(n1383), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[142]) );
  DFFSR \current_reg[150]  ( .D(n1381), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[150]) );
  DFFSR \current_reg[158]  ( .D(n1379), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[158]) );
  DFFSR \current_reg[166]  ( .D(n1377), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[166]) );
  DFFSR \current_reg[174]  ( .D(n1375), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[174]) );
  DFFSR \current_reg[182]  ( .D(n1373), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[182]) );
  DFFSR \current_reg[190]  ( .D(n1371), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[190]) );
  DFFSR \current_reg[198]  ( .D(n1369), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[198]) );
  DFFSR \current_reg[206]  ( .D(n1367), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[206]) );
  DFFSR \current_reg[214]  ( .D(n1365), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[214]) );
  DFFSR \current_reg[222]  ( .D(n1363), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[222]) );
  DFFSR \current_reg[230]  ( .D(n1361), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[230]) );
  DFFSR \current_reg[238]  ( .D(n1359), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[238]) );
  DFFSR \current_reg[246]  ( .D(n1357), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[246]) );
  DFFSR \current_reg[254]  ( .D(n1355), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[254]) );
  DFFSR \current_reg[262]  ( .D(n1353), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[262]) );
  DFFSR \current_reg[270]  ( .D(n1351), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[270]) );
  DFFSR \current_reg[278]  ( .D(n1349), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[278]) );
  DFFSR \current_reg[286]  ( .D(n1347), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[286]) );
  DFFSR \current_reg[294]  ( .D(n1345), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[294]) );
  DFFSR \current_reg[302]  ( .D(n1343), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[302]) );
  DFFSR \current_reg[310]  ( .D(n1341), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[310]) );
  DFFSR \current_reg[318]  ( .D(n1339), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[318]) );
  DFFSR \current_reg[326]  ( .D(n1337), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[326]) );
  DFFSR \current_reg[334]  ( .D(n1335), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[334]) );
  DFFSR \current_reg[342]  ( .D(n1333), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[342]) );
  DFFSR \current_reg[350]  ( .D(n1331), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[350]) );
  DFFSR \current_reg[358]  ( .D(n1329), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[358]) );
  DFFSR \current_reg[366]  ( .D(n1327), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[366]) );
  DFFSR \current_reg[374]  ( .D(n1325), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[374]) );
  DFFSR \current_reg[382]  ( .D(n1323), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[382]) );
  DFFSR \current_reg[390]  ( .D(n1321), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[390]) );
  DFFSR \current_reg[398]  ( .D(n1319), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[398]) );
  DFFSR \current_reg[406]  ( .D(n1317), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[406]) );
  DFFSR \current_reg[414]  ( .D(n1315), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[414]) );
  DFFSR \current_reg[422]  ( .D(n1313), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[422]) );
  DFFSR \current_reg[430]  ( .D(n1311), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[430]) );
  DFFSR \current_reg[438]  ( .D(n1309), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[438]) );
  DFFSR \current_reg[446]  ( .D(n1307), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[446]) );
  DFFSR \current_reg[454]  ( .D(n1305), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[454]) );
  DFFSR \current_reg[462]  ( .D(n1303), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[462]) );
  DFFSR \current_reg[470]  ( .D(n1301), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[470]) );
  DFFSR \current_reg[478]  ( .D(n1299), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[478]) );
  DFFSR \current_reg[486]  ( .D(n1297), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[486]) );
  DFFSR \current_reg[494]  ( .D(n1295), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[494]) );
  DFFSR \current_reg[502]  ( .D(n1293), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[502]) );
  DFFSR \current_reg[510]  ( .D(n1291), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[510]) );
  DFFSR \current_reg[5]  ( .D(n1289), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[5]) );
  DFFSR \current_reg[13]  ( .D(n1287), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[13]) );
  DFFSR \current_reg[21]  ( .D(n1285), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[21]) );
  DFFSR \current_reg[29]  ( .D(n1283), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[29]) );
  DFFSR \current_reg[37]  ( .D(n1281), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[37]) );
  DFFSR \current_reg[45]  ( .D(n1279), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[45]) );
  DFFSR \current_reg[53]  ( .D(n1277), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[53]) );
  DFFSR \current_reg[61]  ( .D(n1275), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[61]) );
  DFFSR \current_reg[69]  ( .D(n1273), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[69]) );
  DFFSR \current_reg[77]  ( .D(n1271), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[77]) );
  DFFSR \current_reg[85]  ( .D(n1269), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[85]) );
  DFFSR \current_reg[93]  ( .D(n1267), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[93]) );
  DFFSR \current_reg[101]  ( .D(n1265), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[101]) );
  DFFSR \current_reg[109]  ( .D(n1263), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[109]) );
  DFFSR \current_reg[117]  ( .D(n1261), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[117]) );
  DFFSR \current_reg[125]  ( .D(n1259), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[125]) );
  DFFSR \current_reg[133]  ( .D(n1257), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[133]) );
  DFFSR \current_reg[141]  ( .D(n1255), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[141]) );
  DFFSR \current_reg[149]  ( .D(n1253), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[149]) );
  DFFSR \current_reg[157]  ( .D(n1251), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[157]) );
  DFFSR \current_reg[165]  ( .D(n1249), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[165]) );
  DFFSR \current_reg[173]  ( .D(n1247), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[173]) );
  DFFSR \current_reg[181]  ( .D(n1245), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[181]) );
  DFFSR \current_reg[189]  ( .D(n1243), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[189]) );
  DFFSR \current_reg[197]  ( .D(n1241), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[197]) );
  DFFSR \current_reg[205]  ( .D(n1239), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[205]) );
  DFFSR \current_reg[213]  ( .D(n1237), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[213]) );
  DFFSR \current_reg[221]  ( .D(n1235), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[221]) );
  DFFSR \current_reg[229]  ( .D(n1233), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[229]) );
  DFFSR \current_reg[237]  ( .D(n1231), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[237]) );
  DFFSR \current_reg[245]  ( .D(n1229), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[245]) );
  DFFSR \current_reg[253]  ( .D(n1227), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[253]) );
  DFFSR \current_reg[261]  ( .D(n1225), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[261]) );
  DFFSR \current_reg[269]  ( .D(n1223), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[269]) );
  DFFSR \current_reg[277]  ( .D(n1221), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[277]) );
  DFFSR \current_reg[285]  ( .D(n1219), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[285]) );
  DFFSR \current_reg[293]  ( .D(n1217), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[293]) );
  DFFSR \current_reg[301]  ( .D(n1215), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[301]) );
  DFFSR \current_reg[309]  ( .D(n1213), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[309]) );
  DFFSR \current_reg[317]  ( .D(n1211), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[317]) );
  DFFSR \current_reg[325]  ( .D(n1209), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[325]) );
  DFFSR \current_reg[333]  ( .D(n1207), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[333]) );
  DFFSR \current_reg[341]  ( .D(n1205), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[341]) );
  DFFSR \current_reg[349]  ( .D(n1203), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[349]) );
  DFFSR \current_reg[357]  ( .D(n1201), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[357]) );
  DFFSR \current_reg[365]  ( .D(n1199), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[365]) );
  DFFSR \current_reg[373]  ( .D(n1197), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[373]) );
  DFFSR \current_reg[381]  ( .D(n1195), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[381]) );
  DFFSR \current_reg[389]  ( .D(n1193), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[389]) );
  DFFSR \current_reg[397]  ( .D(n1191), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[397]) );
  DFFSR \current_reg[405]  ( .D(n1189), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[405]) );
  DFFSR \current_reg[413]  ( .D(n1187), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[413]) );
  DFFSR \current_reg[421]  ( .D(n1185), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[421]) );
  DFFSR \current_reg[429]  ( .D(n1183), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[429]) );
  DFFSR \current_reg[437]  ( .D(n1181), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[437]) );
  DFFSR \current_reg[445]  ( .D(n1179), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[445]) );
  DFFSR \current_reg[453]  ( .D(n1177), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[453]) );
  DFFSR \current_reg[461]  ( .D(n1175), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[461]) );
  DFFSR \current_reg[469]  ( .D(n1173), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[469]) );
  DFFSR \current_reg[477]  ( .D(n1171), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[477]) );
  DFFSR \current_reg[485]  ( .D(n1169), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[485]) );
  DFFSR \current_reg[493]  ( .D(n1167), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[493]) );
  DFFSR \current_reg[501]  ( .D(n1165), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[501]) );
  DFFSR \current_reg[509]  ( .D(n1163), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[509]) );
  DFFSR \current_reg[4]  ( .D(n1161), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[4]) );
  DFFSR \current_reg[12]  ( .D(n1159), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[12]) );
  DFFSR \current_reg[20]  ( .D(n1157), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[20]) );
  DFFSR \current_reg[28]  ( .D(n1155), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[28]) );
  DFFSR \current_reg[36]  ( .D(n1153), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[36]) );
  DFFSR \current_reg[44]  ( .D(n1151), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[44]) );
  DFFSR \current_reg[52]  ( .D(n1149), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[52]) );
  DFFSR \current_reg[60]  ( .D(n1147), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[60]) );
  DFFSR \current_reg[68]  ( .D(n1145), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[68]) );
  DFFSR \current_reg[76]  ( .D(n1143), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[76]) );
  DFFSR \current_reg[84]  ( .D(n1141), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[84]) );
  DFFSR \current_reg[92]  ( .D(n1139), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[92]) );
  DFFSR \current_reg[100]  ( .D(n1137), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[100]) );
  DFFSR \current_reg[108]  ( .D(n1135), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[108]) );
  DFFSR \current_reg[116]  ( .D(n1133), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[116]) );
  DFFSR \current_reg[124]  ( .D(n1131), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[124]) );
  DFFSR \current_reg[132]  ( .D(n1129), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[132]) );
  DFFSR \current_reg[140]  ( .D(n1127), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[140]) );
  DFFSR \current_reg[148]  ( .D(n1125), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[148]) );
  DFFSR \current_reg[156]  ( .D(n1123), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[156]) );
  DFFSR \current_reg[164]  ( .D(n1121), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[164]) );
  DFFSR \current_reg[172]  ( .D(n1119), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[172]) );
  DFFSR \current_reg[180]  ( .D(n1117), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[180]) );
  DFFSR \current_reg[188]  ( .D(n1115), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[188]) );
  DFFSR \current_reg[196]  ( .D(n1113), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[196]) );
  DFFSR \current_reg[204]  ( .D(n1111), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[204]) );
  DFFSR \current_reg[212]  ( .D(n1109), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[212]) );
  DFFSR \current_reg[220]  ( .D(n1107), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[220]) );
  DFFSR \current_reg[228]  ( .D(n1105), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[228]) );
  DFFSR \current_reg[236]  ( .D(n1103), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[236]) );
  DFFSR \current_reg[244]  ( .D(n1101), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[244]) );
  DFFSR \current_reg[252]  ( .D(n1099), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[252]) );
  DFFSR \current_reg[260]  ( .D(n1097), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[260]) );
  DFFSR \current_reg[268]  ( .D(n1095), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[268]) );
  DFFSR \current_reg[276]  ( .D(n1093), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[276]) );
  DFFSR \current_reg[284]  ( .D(n1091), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[284]) );
  DFFSR \current_reg[292]  ( .D(n1089), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[292]) );
  DFFSR \current_reg[300]  ( .D(n1087), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[300]) );
  DFFSR \current_reg[308]  ( .D(n1085), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[308]) );
  DFFSR \current_reg[316]  ( .D(n1083), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[316]) );
  DFFSR \current_reg[324]  ( .D(n1081), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[324]) );
  DFFSR \current_reg[332]  ( .D(n1079), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[332]) );
  DFFSR \current_reg[340]  ( .D(n1077), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[340]) );
  DFFSR \current_reg[348]  ( .D(n1075), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[348]) );
  DFFSR \current_reg[356]  ( .D(n1073), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[356]) );
  DFFSR \current_reg[364]  ( .D(n1071), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[364]) );
  DFFSR \current_reg[372]  ( .D(n1069), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[372]) );
  DFFSR \current_reg[380]  ( .D(n1067), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[380]) );
  DFFSR \current_reg[388]  ( .D(n1065), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[388]) );
  DFFSR \current_reg[396]  ( .D(n1063), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[396]) );
  DFFSR \current_reg[404]  ( .D(n1061), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[404]) );
  DFFSR \current_reg[412]  ( .D(n1059), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[412]) );
  DFFSR \current_reg[420]  ( .D(n1057), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[420]) );
  DFFSR \current_reg[428]  ( .D(n1055), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[428]) );
  DFFSR \current_reg[436]  ( .D(n1053), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[436]) );
  DFFSR \current_reg[444]  ( .D(n1051), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[444]) );
  DFFSR \current_reg[452]  ( .D(n1049), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[452]) );
  DFFSR \current_reg[460]  ( .D(n1047), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[460]) );
  DFFSR \current_reg[468]  ( .D(n1045), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[468]) );
  DFFSR \current_reg[476]  ( .D(n1043), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[476]) );
  DFFSR \current_reg[484]  ( .D(n1041), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[484]) );
  DFFSR \current_reg[492]  ( .D(n1039), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[492]) );
  DFFSR \current_reg[500]  ( .D(n1037), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[500]) );
  DFFSR \current_reg[508]  ( .D(n1035), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[508]) );
  DFFSR \current_reg[3]  ( .D(n1033), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[3]) );
  DFFSR \current_reg[11]  ( .D(n1031), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[11]) );
  DFFSR \current_reg[19]  ( .D(n1029), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[19]) );
  DFFSR \current_reg[27]  ( .D(n1027), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[27]) );
  DFFSR \current_reg[35]  ( .D(n1025), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[35]) );
  DFFSR \current_reg[43]  ( .D(n1023), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[43]) );
  DFFSR \current_reg[51]  ( .D(n1021), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[51]) );
  DFFSR \current_reg[59]  ( .D(n1019), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[59]) );
  DFFSR \current_reg[67]  ( .D(n1017), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[67]) );
  DFFSR \current_reg[75]  ( .D(n1015), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[75]) );
  DFFSR \current_reg[83]  ( .D(n1013), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[83]) );
  DFFSR \current_reg[91]  ( .D(n1011), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[91]) );
  DFFSR \current_reg[99]  ( .D(n1009), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[99]) );
  DFFSR \current_reg[107]  ( .D(n1007), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[107]) );
  DFFSR \current_reg[115]  ( .D(n1005), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[115]) );
  DFFSR \current_reg[123]  ( .D(n1003), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[123]) );
  DFFSR \current_reg[131]  ( .D(n1001), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[131]) );
  DFFSR \current_reg[139]  ( .D(n999), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[139]) );
  DFFSR \current_reg[147]  ( .D(n997), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[147]) );
  DFFSR \current_reg[155]  ( .D(n995), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[155]) );
  DFFSR \current_reg[163]  ( .D(n993), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[163]) );
  DFFSR \current_reg[171]  ( .D(n991), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[171]) );
  DFFSR \current_reg[179]  ( .D(n989), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[179]) );
  DFFSR \current_reg[187]  ( .D(n987), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[187]) );
  DFFSR \current_reg[195]  ( .D(n985), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[195]) );
  DFFSR \current_reg[203]  ( .D(n983), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[203]) );
  DFFSR \current_reg[211]  ( .D(n981), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[211]) );
  DFFSR \current_reg[219]  ( .D(n979), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[219]) );
  DFFSR \current_reg[227]  ( .D(n977), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[227]) );
  DFFSR \current_reg[235]  ( .D(n975), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[235]) );
  DFFSR \current_reg[243]  ( .D(n973), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[243]) );
  DFFSR \current_reg[251]  ( .D(n971), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[251]) );
  DFFSR \current_reg[259]  ( .D(n969), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[259]) );
  DFFSR \current_reg[267]  ( .D(n967), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[267]) );
  DFFSR \current_reg[275]  ( .D(n965), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[275]) );
  DFFSR \current_reg[283]  ( .D(n963), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[283]) );
  DFFSR \current_reg[291]  ( .D(n961), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[291]) );
  DFFSR \current_reg[299]  ( .D(n959), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[299]) );
  DFFSR \current_reg[307]  ( .D(n957), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[307]) );
  DFFSR \current_reg[315]  ( .D(n955), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[315]) );
  DFFSR \current_reg[323]  ( .D(n953), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[323]) );
  DFFSR \current_reg[331]  ( .D(n951), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[331]) );
  DFFSR \current_reg[339]  ( .D(n949), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[339]) );
  DFFSR \current_reg[347]  ( .D(n947), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[347]) );
  DFFSR \current_reg[355]  ( .D(n945), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[355]) );
  DFFSR \current_reg[363]  ( .D(n943), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[363]) );
  DFFSR \current_reg[371]  ( .D(n941), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[371]) );
  DFFSR \current_reg[379]  ( .D(n939), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[379]) );
  DFFSR \current_reg[387]  ( .D(n937), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[387]) );
  DFFSR \current_reg[395]  ( .D(n935), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[395]) );
  DFFSR \current_reg[403]  ( .D(n933), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[403]) );
  DFFSR \current_reg[411]  ( .D(n931), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[411]) );
  DFFSR \current_reg[419]  ( .D(n929), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[419]) );
  DFFSR \current_reg[427]  ( .D(n927), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[427]) );
  DFFSR \current_reg[435]  ( .D(n925), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[435]) );
  DFFSR \current_reg[443]  ( .D(n923), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[443]) );
  DFFSR \current_reg[451]  ( .D(n921), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[451]) );
  DFFSR \current_reg[459]  ( .D(n919), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[459]) );
  DFFSR \current_reg[467]  ( .D(n917), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[467]) );
  DFFSR \current_reg[475]  ( .D(n915), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[475]) );
  DFFSR \current_reg[483]  ( .D(n913), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[483]) );
  DFFSR \current_reg[491]  ( .D(n911), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[491]) );
  DFFSR \current_reg[499]  ( .D(n909), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[499]) );
  DFFSR \current_reg[507]  ( .D(n907), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[507]) );
  DFFSR \current_reg[2]  ( .D(n905), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[2]) );
  DFFSR \current_reg[10]  ( .D(n903), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[10]) );
  DFFSR \current_reg[18]  ( .D(n901), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[18]) );
  DFFSR \current_reg[26]  ( .D(n899), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[26]) );
  DFFSR \current_reg[34]  ( .D(n897), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[34]) );
  DFFSR \current_reg[42]  ( .D(n895), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[42]) );
  DFFSR \current_reg[50]  ( .D(n893), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[50]) );
  DFFSR \current_reg[58]  ( .D(n891), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[58]) );
  DFFSR \current_reg[66]  ( .D(n889), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[66]) );
  DFFSR \current_reg[74]  ( .D(n887), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[74]) );
  DFFSR \current_reg[82]  ( .D(n885), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[82]) );
  DFFSR \current_reg[90]  ( .D(n883), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[90]) );
  DFFSR \current_reg[98]  ( .D(n881), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[98]) );
  DFFSR \current_reg[106]  ( .D(n879), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[106]) );
  DFFSR \current_reg[114]  ( .D(n877), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[114]) );
  DFFSR \current_reg[122]  ( .D(n875), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[122]) );
  DFFSR \current_reg[130]  ( .D(n873), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[130]) );
  DFFSR \current_reg[138]  ( .D(n871), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[138]) );
  DFFSR \current_reg[146]  ( .D(n869), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[146]) );
  DFFSR \current_reg[154]  ( .D(n867), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[154]) );
  DFFSR \current_reg[162]  ( .D(n865), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[162]) );
  DFFSR \current_reg[170]  ( .D(n863), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[170]) );
  DFFSR \current_reg[178]  ( .D(n861), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[178]) );
  DFFSR \current_reg[186]  ( .D(n859), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[186]) );
  DFFSR \current_reg[194]  ( .D(n857), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[194]) );
  DFFSR \current_reg[202]  ( .D(n855), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[202]) );
  DFFSR \current_reg[210]  ( .D(n853), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[210]) );
  DFFSR \current_reg[218]  ( .D(n851), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[218]) );
  DFFSR \current_reg[226]  ( .D(n849), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[226]) );
  DFFSR \current_reg[234]  ( .D(n847), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[234]) );
  DFFSR \current_reg[242]  ( .D(n845), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[242]) );
  DFFSR \current_reg[250]  ( .D(n843), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[250]) );
  DFFSR \current_reg[258]  ( .D(n841), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[258]) );
  DFFSR \current_reg[266]  ( .D(n839), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[266]) );
  DFFSR \current_reg[274]  ( .D(n837), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[274]) );
  DFFSR \current_reg[282]  ( .D(n835), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[282]) );
  DFFSR \current_reg[290]  ( .D(n833), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[290]) );
  DFFSR \current_reg[298]  ( .D(n831), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[298]) );
  DFFSR \current_reg[306]  ( .D(n829), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[306]) );
  DFFSR \current_reg[314]  ( .D(n827), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[314]) );
  DFFSR \current_reg[322]  ( .D(n825), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[322]) );
  DFFSR \current_reg[330]  ( .D(n823), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[330]) );
  DFFSR \current_reg[338]  ( .D(n821), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[338]) );
  DFFSR \current_reg[346]  ( .D(n819), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[346]) );
  DFFSR \current_reg[354]  ( .D(n817), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[354]) );
  DFFSR \current_reg[362]  ( .D(n815), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[362]) );
  DFFSR \current_reg[370]  ( .D(n813), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[370]) );
  DFFSR \current_reg[378]  ( .D(n811), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[378]) );
  DFFSR \current_reg[386]  ( .D(n809), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[386]) );
  DFFSR \current_reg[394]  ( .D(n807), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[394]) );
  DFFSR \current_reg[402]  ( .D(n805), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[402]) );
  DFFSR \current_reg[410]  ( .D(n803), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[410]) );
  DFFSR \current_reg[418]  ( .D(n801), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[418]) );
  DFFSR \current_reg[426]  ( .D(n799), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[426]) );
  DFFSR \current_reg[434]  ( .D(n797), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[434]) );
  DFFSR \current_reg[442]  ( .D(n795), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[442]) );
  DFFSR \current_reg[450]  ( .D(n793), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[450]) );
  DFFSR \current_reg[458]  ( .D(n791), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[458]) );
  DFFSR \current_reg[466]  ( .D(n789), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[466]) );
  DFFSR \current_reg[474]  ( .D(n787), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[474]) );
  DFFSR \current_reg[482]  ( .D(n785), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[482]) );
  DFFSR \current_reg[490]  ( .D(n783), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[490]) );
  DFFSR \current_reg[498]  ( .D(n781), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[498]) );
  DFFSR \current_reg[506]  ( .D(n779), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[506]) );
  DFFSR \current_reg[1]  ( .D(n777), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[1]) );
  DFFSR \current_reg[9]  ( .D(n775), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[9]) );
  DFFSR \current_reg[17]  ( .D(n773), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[17]) );
  DFFSR \current_reg[25]  ( .D(n771), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[25]) );
  DFFSR \current_reg[33]  ( .D(n769), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[33]) );
  DFFSR \current_reg[41]  ( .D(n767), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[41]) );
  DFFSR \current_reg[49]  ( .D(n765), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[49]) );
  DFFSR \current_reg[57]  ( .D(n763), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[57]) );
  DFFSR \current_reg[65]  ( .D(n761), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[65]) );
  DFFSR \current_reg[73]  ( .D(n759), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[73]) );
  DFFSR \current_reg[81]  ( .D(n757), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[81]) );
  DFFSR \current_reg[89]  ( .D(n755), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[89]) );
  DFFSR \current_reg[97]  ( .D(n753), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[97]) );
  DFFSR \current_reg[105]  ( .D(n751), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[105]) );
  DFFSR \current_reg[113]  ( .D(n749), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[113]) );
  DFFSR \current_reg[121]  ( .D(n747), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[121]) );
  DFFSR \current_reg[129]  ( .D(n745), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[129]) );
  DFFSR \current_reg[137]  ( .D(n743), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[137]) );
  DFFSR \current_reg[145]  ( .D(n741), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[145]) );
  DFFSR \current_reg[153]  ( .D(n739), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[153]) );
  DFFSR \current_reg[161]  ( .D(n737), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[161]) );
  DFFSR \current_reg[169]  ( .D(n735), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[169]) );
  DFFSR \current_reg[177]  ( .D(n733), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[177]) );
  DFFSR \current_reg[185]  ( .D(n731), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[185]) );
  DFFSR \current_reg[193]  ( .D(n729), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[193]) );
  DFFSR \current_reg[201]  ( .D(n727), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[201]) );
  DFFSR \current_reg[209]  ( .D(n725), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[209]) );
  DFFSR \current_reg[217]  ( .D(n723), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[217]) );
  DFFSR \current_reg[225]  ( .D(n721), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[225]) );
  DFFSR \current_reg[233]  ( .D(n719), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[233]) );
  DFFSR \current_reg[241]  ( .D(n717), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[241]) );
  DFFSR \current_reg[249]  ( .D(n715), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[249]) );
  DFFSR \current_reg[257]  ( .D(n713), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[257]) );
  DFFSR \current_reg[265]  ( .D(n711), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[265]) );
  DFFSR \current_reg[273]  ( .D(n709), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[273]) );
  DFFSR \current_reg[281]  ( .D(n707), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[281]) );
  DFFSR \current_reg[289]  ( .D(n705), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[289]) );
  DFFSR \current_reg[297]  ( .D(n703), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[297]) );
  DFFSR \current_reg[305]  ( .D(n701), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[305]) );
  DFFSR \current_reg[313]  ( .D(n699), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[313]) );
  DFFSR \current_reg[321]  ( .D(n697), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[321]) );
  DFFSR \current_reg[329]  ( .D(n695), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[329]) );
  DFFSR \current_reg[337]  ( .D(n693), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[337]) );
  DFFSR \current_reg[345]  ( .D(n691), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[345]) );
  DFFSR \current_reg[353]  ( .D(n689), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[353]) );
  DFFSR \current_reg[361]  ( .D(n687), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[361]) );
  DFFSR \current_reg[369]  ( .D(n685), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[369]) );
  DFFSR \current_reg[377]  ( .D(n683), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[377]) );
  DFFSR \current_reg[385]  ( .D(n681), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[385]) );
  DFFSR \current_reg[393]  ( .D(n679), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[393]) );
  DFFSR \current_reg[401]  ( .D(n677), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[401]) );
  DFFSR \current_reg[409]  ( .D(n675), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[409]) );
  DFFSR \current_reg[417]  ( .D(n673), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[417]) );
  DFFSR \current_reg[425]  ( .D(n671), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[425]) );
  DFFSR \current_reg[433]  ( .D(n669), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[433]) );
  DFFSR \current_reg[441]  ( .D(n667), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[441]) );
  DFFSR \current_reg[449]  ( .D(n665), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[449]) );
  DFFSR \current_reg[457]  ( .D(n663), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[457]) );
  DFFSR \current_reg[465]  ( .D(n661), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[465]) );
  DFFSR \current_reg[473]  ( .D(n659), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[473]) );
  DFFSR \current_reg[481]  ( .D(n657), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[481]) );
  DFFSR \current_reg[489]  ( .D(n655), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[489]) );
  DFFSR \current_reg[497]  ( .D(n653), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[497]) );
  DFFSR \current_reg[505]  ( .D(n651), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[505]) );
  DFFSR \current_reg[0]  ( .D(n649), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[0]) );
  DFFSR \current_reg[8]  ( .D(n647), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[8]) );
  DFFSR \current_reg[16]  ( .D(n645), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[16]) );
  DFFSR \current_reg[24]  ( .D(n643), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[24]) );
  DFFSR \current_reg[32]  ( .D(n641), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[32]) );
  DFFSR \current_reg[40]  ( .D(n639), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[40]) );
  DFFSR \current_reg[48]  ( .D(n637), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[48]) );
  DFFSR \current_reg[56]  ( .D(n635), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[56]) );
  DFFSR \current_reg[64]  ( .D(n633), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[64]) );
  DFFSR \current_reg[72]  ( .D(n631), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[72]) );
  DFFSR \current_reg[80]  ( .D(n629), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[80]) );
  DFFSR \current_reg[88]  ( .D(n627), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[88]) );
  DFFSR \current_reg[96]  ( .D(n625), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[96]) );
  DFFSR \current_reg[104]  ( .D(n623), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[104]) );
  DFFSR \current_reg[112]  ( .D(n621), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[112]) );
  DFFSR \current_reg[120]  ( .D(n619), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[120]) );
  DFFSR \current_reg[128]  ( .D(n617), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[128]) );
  DFFSR \current_reg[136]  ( .D(n615), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[136]) );
  DFFSR \current_reg[144]  ( .D(n613), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[144]) );
  DFFSR \current_reg[152]  ( .D(n611), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[152]) );
  DFFSR \current_reg[160]  ( .D(n609), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[160]) );
  DFFSR \current_reg[168]  ( .D(n607), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[168]) );
  DFFSR \current_reg[176]  ( .D(n605), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[176]) );
  DFFSR \current_reg[184]  ( .D(n603), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[184]) );
  DFFSR \current_reg[192]  ( .D(n601), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[192]) );
  DFFSR \current_reg[200]  ( .D(n599), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[200]) );
  DFFSR \current_reg[208]  ( .D(n597), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[208]) );
  DFFSR \current_reg[216]  ( .D(n595), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[216]) );
  DFFSR \current_reg[224]  ( .D(n593), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[224]) );
  DFFSR \current_reg[232]  ( .D(n591), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[232]) );
  DFFSR \current_reg[240]  ( .D(n589), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[240]) );
  DFFSR \current_reg[248]  ( .D(n587), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[248]) );
  DFFSR \current_reg[256]  ( .D(n585), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[256]) );
  DFFSR \current_reg[264]  ( .D(n583), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[264]) );
  DFFSR \current_reg[272]  ( .D(n581), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[272]) );
  DFFSR \current_reg[280]  ( .D(n579), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[280]) );
  DFFSR \current_reg[288]  ( .D(n577), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[288]) );
  DFFSR \current_reg[296]  ( .D(n575), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[296]) );
  DFFSR \current_reg[304]  ( .D(n573), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[304]) );
  DFFSR \current_reg[312]  ( .D(n571), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[312]) );
  DFFSR \current_reg[320]  ( .D(n569), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[320]) );
  DFFSR \current_reg[328]  ( .D(n567), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[328]) );
  DFFSR \current_reg[336]  ( .D(n565), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[336]) );
  DFFSR \current_reg[344]  ( .D(n563), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[344]) );
  DFFSR \current_reg[352]  ( .D(n561), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[352]) );
  DFFSR \current_reg[360]  ( .D(n559), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[360]) );
  DFFSR \current_reg[368]  ( .D(n557), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[368]) );
  DFFSR \current_reg[376]  ( .D(n555), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[376]) );
  DFFSR \current_reg[384]  ( .D(n553), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[384]) );
  DFFSR \current_reg[392]  ( .D(n551), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[392]) );
  DFFSR \current_reg[400]  ( .D(n549), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[400]) );
  DFFSR \current_reg[408]  ( .D(n547), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[408]) );
  DFFSR \current_reg[416]  ( .D(n545), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[416]) );
  DFFSR \current_reg[424]  ( .D(n543), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[424]) );
  DFFSR \current_reg[432]  ( .D(n541), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[432]) );
  DFFSR \current_reg[440]  ( .D(n539), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[440]) );
  DFFSR \current_reg[448]  ( .D(n537), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[448]) );
  DFFSR \current_reg[456]  ( .D(n535), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[456]) );
  DFFSR \current_reg[464]  ( .D(n533), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[464]) );
  DFFSR \current_reg[472]  ( .D(n531), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[472]) );
  DFFSR \current_reg[480]  ( .D(n529), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[480]) );
  DFFSR \current_reg[488]  ( .D(n527), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[488]) );
  DFFSR \current_reg[496]  ( .D(n525), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[496]) );
  DFFSR \current_reg[504]  ( .D(n523), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        data_out[504]) );
  INVX1 U1547 ( .A(n1546), .Y(n999) );
  MUX2X1 U1548 ( .B(data_out[139]), .A(data_out[131]), .S(shift_en), .Y(n1546)
         );
  INVX1 U1549 ( .A(n1547), .Y(n997) );
  MUX2X1 U1550 ( .B(data_out[147]), .A(data_out[139]), .S(shift_en), .Y(n1547)
         );
  INVX1 U1551 ( .A(n1548), .Y(n995) );
  MUX2X1 U1552 ( .B(data_out[155]), .A(data_out[147]), .S(shift_en), .Y(n1548)
         );
  INVX1 U1553 ( .A(n1549), .Y(n993) );
  MUX2X1 U1554 ( .B(data_out[163]), .A(data_out[155]), .S(shift_en), .Y(n1549)
         );
  INVX1 U1555 ( .A(n1550), .Y(n991) );
  MUX2X1 U1556 ( .B(data_out[171]), .A(data_out[163]), .S(shift_en), .Y(n1550)
         );
  INVX1 U1557 ( .A(n1551), .Y(n989) );
  MUX2X1 U1558 ( .B(data_out[179]), .A(data_out[171]), .S(shift_en), .Y(n1551)
         );
  INVX1 U1559 ( .A(n1552), .Y(n987) );
  MUX2X1 U1560 ( .B(data_out[187]), .A(data_out[179]), .S(shift_en), .Y(n1552)
         );
  INVX1 U1561 ( .A(n1553), .Y(n985) );
  MUX2X1 U1562 ( .B(data_out[195]), .A(data_out[187]), .S(shift_en), .Y(n1553)
         );
  INVX1 U1563 ( .A(n1554), .Y(n983) );
  MUX2X1 U1564 ( .B(data_out[203]), .A(data_out[195]), .S(shift_en), .Y(n1554)
         );
  INVX1 U1565 ( .A(n1555), .Y(n981) );
  MUX2X1 U1566 ( .B(data_out[211]), .A(data_out[203]), .S(shift_en), .Y(n1555)
         );
  INVX1 U1567 ( .A(n1556), .Y(n979) );
  MUX2X1 U1568 ( .B(data_out[219]), .A(data_out[211]), .S(shift_en), .Y(n1556)
         );
  INVX1 U1569 ( .A(n1557), .Y(n977) );
  MUX2X1 U1570 ( .B(data_out[227]), .A(data_out[219]), .S(shift_en), .Y(n1557)
         );
  INVX1 U1571 ( .A(n1558), .Y(n975) );
  MUX2X1 U1572 ( .B(data_out[235]), .A(data_out[227]), .S(shift_en), .Y(n1558)
         );
  INVX1 U1573 ( .A(n1559), .Y(n973) );
  MUX2X1 U1574 ( .B(data_out[243]), .A(data_out[235]), .S(shift_en), .Y(n1559)
         );
  INVX1 U1575 ( .A(n1560), .Y(n971) );
  MUX2X1 U1576 ( .B(data_out[251]), .A(data_out[243]), .S(shift_en), .Y(n1560)
         );
  INVX1 U1577 ( .A(n1561), .Y(n969) );
  MUX2X1 U1578 ( .B(data_out[259]), .A(data_out[251]), .S(shift_en), .Y(n1561)
         );
  INVX1 U1579 ( .A(n1562), .Y(n967) );
  MUX2X1 U1580 ( .B(data_out[267]), .A(data_out[259]), .S(shift_en), .Y(n1562)
         );
  INVX1 U1581 ( .A(n1563), .Y(n965) );
  MUX2X1 U1582 ( .B(data_out[275]), .A(data_out[267]), .S(shift_en), .Y(n1563)
         );
  INVX1 U1583 ( .A(n1564), .Y(n963) );
  MUX2X1 U1584 ( .B(data_out[283]), .A(data_out[275]), .S(shift_en), .Y(n1564)
         );
  INVX1 U1585 ( .A(n1565), .Y(n961) );
  MUX2X1 U1586 ( .B(data_out[291]), .A(data_out[283]), .S(shift_en), .Y(n1565)
         );
  INVX1 U1587 ( .A(n1566), .Y(n959) );
  MUX2X1 U1588 ( .B(data_out[299]), .A(data_out[291]), .S(shift_en), .Y(n1566)
         );
  INVX1 U1589 ( .A(n1567), .Y(n957) );
  MUX2X1 U1590 ( .B(data_out[307]), .A(data_out[299]), .S(shift_en), .Y(n1567)
         );
  INVX1 U1591 ( .A(n1568), .Y(n955) );
  MUX2X1 U1592 ( .B(data_out[315]), .A(data_out[307]), .S(shift_en), .Y(n1568)
         );
  INVX1 U1593 ( .A(n1569), .Y(n953) );
  MUX2X1 U1594 ( .B(data_out[323]), .A(data_out[315]), .S(shift_en), .Y(n1569)
         );
  INVX1 U1595 ( .A(n1570), .Y(n951) );
  MUX2X1 U1596 ( .B(data_out[331]), .A(data_out[323]), .S(shift_en), .Y(n1570)
         );
  INVX1 U1597 ( .A(n1571), .Y(n949) );
  MUX2X1 U1598 ( .B(data_out[339]), .A(data_out[331]), .S(shift_en), .Y(n1571)
         );
  INVX1 U1599 ( .A(n1572), .Y(n947) );
  MUX2X1 U1600 ( .B(data_out[347]), .A(data_out[339]), .S(shift_en), .Y(n1572)
         );
  INVX1 U1601 ( .A(n1573), .Y(n945) );
  MUX2X1 U1602 ( .B(data_out[355]), .A(data_out[347]), .S(shift_en), .Y(n1573)
         );
  INVX1 U1603 ( .A(n1574), .Y(n943) );
  MUX2X1 U1604 ( .B(data_out[363]), .A(data_out[355]), .S(shift_en), .Y(n1574)
         );
  INVX1 U1605 ( .A(n1575), .Y(n941) );
  MUX2X1 U1606 ( .B(data_out[371]), .A(data_out[363]), .S(shift_en), .Y(n1575)
         );
  INVX1 U1607 ( .A(n1576), .Y(n939) );
  MUX2X1 U1608 ( .B(data_out[379]), .A(data_out[371]), .S(shift_en), .Y(n1576)
         );
  INVX1 U1609 ( .A(n1577), .Y(n937) );
  MUX2X1 U1610 ( .B(data_out[387]), .A(data_out[379]), .S(shift_en), .Y(n1577)
         );
  INVX1 U1611 ( .A(n1578), .Y(n935) );
  MUX2X1 U1612 ( .B(data_out[395]), .A(data_out[387]), .S(shift_en), .Y(n1578)
         );
  INVX1 U1613 ( .A(n1579), .Y(n933) );
  MUX2X1 U1614 ( .B(data_out[403]), .A(data_out[395]), .S(shift_en), .Y(n1579)
         );
  INVX1 U1615 ( .A(n1580), .Y(n931) );
  MUX2X1 U1616 ( .B(data_out[411]), .A(data_out[403]), .S(shift_en), .Y(n1580)
         );
  INVX1 U1617 ( .A(n1581), .Y(n929) );
  MUX2X1 U1618 ( .B(data_out[419]), .A(data_out[411]), .S(shift_en), .Y(n1581)
         );
  INVX1 U1619 ( .A(n1582), .Y(n927) );
  MUX2X1 U1620 ( .B(data_out[427]), .A(data_out[419]), .S(shift_en), .Y(n1582)
         );
  INVX1 U1621 ( .A(n1583), .Y(n925) );
  MUX2X1 U1622 ( .B(data_out[435]), .A(data_out[427]), .S(shift_en), .Y(n1583)
         );
  INVX1 U1623 ( .A(n1584), .Y(n923) );
  MUX2X1 U1624 ( .B(data_out[443]), .A(data_out[435]), .S(shift_en), .Y(n1584)
         );
  INVX1 U1625 ( .A(n1585), .Y(n921) );
  MUX2X1 U1626 ( .B(data_out[451]), .A(data_out[443]), .S(shift_en), .Y(n1585)
         );
  INVX1 U1627 ( .A(n1586), .Y(n919) );
  MUX2X1 U1628 ( .B(data_out[459]), .A(data_out[451]), .S(shift_en), .Y(n1586)
         );
  INVX1 U1629 ( .A(n1587), .Y(n917) );
  MUX2X1 U1630 ( .B(data_out[467]), .A(data_out[459]), .S(shift_en), .Y(n1587)
         );
  INVX1 U1631 ( .A(n1588), .Y(n915) );
  MUX2X1 U1632 ( .B(data_out[475]), .A(data_out[467]), .S(shift_en), .Y(n1588)
         );
  INVX1 U1633 ( .A(n1589), .Y(n913) );
  MUX2X1 U1634 ( .B(data_out[483]), .A(data_out[475]), .S(shift_en), .Y(n1589)
         );
  INVX1 U1635 ( .A(n1590), .Y(n911) );
  MUX2X1 U1636 ( .B(data_out[491]), .A(data_out[483]), .S(shift_en), .Y(n1590)
         );
  INVX1 U1637 ( .A(n1591), .Y(n909) );
  MUX2X1 U1638 ( .B(data_out[499]), .A(data_out[491]), .S(shift_en), .Y(n1591)
         );
  INVX1 U1639 ( .A(n1592), .Y(n907) );
  MUX2X1 U1640 ( .B(data_out[507]), .A(data_out[499]), .S(shift_en), .Y(n1592)
         );
  INVX1 U1641 ( .A(n1593), .Y(n905) );
  MUX2X1 U1642 ( .B(data_out[2]), .A(data_in[2]), .S(shift_en), .Y(n1593) );
  INVX1 U1643 ( .A(n1594), .Y(n903) );
  MUX2X1 U1644 ( .B(data_out[10]), .A(data_out[2]), .S(shift_en), .Y(n1594) );
  INVX1 U1645 ( .A(n1595), .Y(n901) );
  MUX2X1 U1646 ( .B(data_out[18]), .A(data_out[10]), .S(shift_en), .Y(n1595)
         );
  INVX1 U1647 ( .A(n1596), .Y(n899) );
  MUX2X1 U1648 ( .B(data_out[26]), .A(data_out[18]), .S(shift_en), .Y(n1596)
         );
  INVX1 U1649 ( .A(n1597), .Y(n897) );
  MUX2X1 U1650 ( .B(data_out[34]), .A(data_out[26]), .S(shift_en), .Y(n1597)
         );
  INVX1 U1651 ( .A(n1598), .Y(n895) );
  MUX2X1 U1652 ( .B(data_out[42]), .A(data_out[34]), .S(shift_en), .Y(n1598)
         );
  INVX1 U1653 ( .A(n1599), .Y(n893) );
  MUX2X1 U1654 ( .B(data_out[50]), .A(data_out[42]), .S(shift_en), .Y(n1599)
         );
  INVX1 U1655 ( .A(n1600), .Y(n891) );
  MUX2X1 U1656 ( .B(data_out[58]), .A(data_out[50]), .S(shift_en), .Y(n1600)
         );
  INVX1 U1657 ( .A(n1601), .Y(n889) );
  MUX2X1 U1658 ( .B(data_out[66]), .A(data_out[58]), .S(shift_en), .Y(n1601)
         );
  INVX1 U1659 ( .A(n1602), .Y(n887) );
  MUX2X1 U1660 ( .B(data_out[74]), .A(data_out[66]), .S(shift_en), .Y(n1602)
         );
  INVX1 U1661 ( .A(n1603), .Y(n885) );
  MUX2X1 U1662 ( .B(data_out[82]), .A(data_out[74]), .S(shift_en), .Y(n1603)
         );
  INVX1 U1663 ( .A(n1604), .Y(n883) );
  MUX2X1 U1664 ( .B(data_out[90]), .A(data_out[82]), .S(shift_en), .Y(n1604)
         );
  INVX1 U1665 ( .A(n1605), .Y(n881) );
  MUX2X1 U1666 ( .B(data_out[98]), .A(data_out[90]), .S(shift_en), .Y(n1605)
         );
  INVX1 U1667 ( .A(n1606), .Y(n879) );
  MUX2X1 U1668 ( .B(data_out[106]), .A(data_out[98]), .S(shift_en), .Y(n1606)
         );
  INVX1 U1669 ( .A(n1607), .Y(n877) );
  MUX2X1 U1670 ( .B(data_out[114]), .A(data_out[106]), .S(shift_en), .Y(n1607)
         );
  INVX1 U1671 ( .A(n1608), .Y(n875) );
  MUX2X1 U1672 ( .B(data_out[122]), .A(data_out[114]), .S(shift_en), .Y(n1608)
         );
  INVX1 U1673 ( .A(n1609), .Y(n873) );
  MUX2X1 U1674 ( .B(data_out[130]), .A(data_out[122]), .S(shift_en), .Y(n1609)
         );
  INVX1 U1675 ( .A(n1610), .Y(n871) );
  MUX2X1 U1676 ( .B(data_out[138]), .A(data_out[130]), .S(shift_en), .Y(n1610)
         );
  INVX1 U1677 ( .A(n1611), .Y(n869) );
  MUX2X1 U1678 ( .B(data_out[146]), .A(data_out[138]), .S(shift_en), .Y(n1611)
         );
  INVX1 U1679 ( .A(n1612), .Y(n867) );
  MUX2X1 U1680 ( .B(data_out[154]), .A(data_out[146]), .S(shift_en), .Y(n1612)
         );
  INVX1 U1681 ( .A(n1613), .Y(n865) );
  MUX2X1 U1682 ( .B(data_out[162]), .A(data_out[154]), .S(shift_en), .Y(n1613)
         );
  INVX1 U1683 ( .A(n1614), .Y(n863) );
  MUX2X1 U1684 ( .B(data_out[170]), .A(data_out[162]), .S(shift_en), .Y(n1614)
         );
  INVX1 U1685 ( .A(n1615), .Y(n861) );
  MUX2X1 U1686 ( .B(data_out[178]), .A(data_out[170]), .S(shift_en), .Y(n1615)
         );
  INVX1 U1687 ( .A(n1616), .Y(n859) );
  MUX2X1 U1688 ( .B(data_out[186]), .A(data_out[178]), .S(shift_en), .Y(n1616)
         );
  INVX1 U1689 ( .A(n1617), .Y(n857) );
  MUX2X1 U1690 ( .B(data_out[194]), .A(data_out[186]), .S(shift_en), .Y(n1617)
         );
  INVX1 U1691 ( .A(n1618), .Y(n855) );
  MUX2X1 U1692 ( .B(data_out[202]), .A(data_out[194]), .S(shift_en), .Y(n1618)
         );
  INVX1 U1693 ( .A(n1619), .Y(n853) );
  MUX2X1 U1694 ( .B(data_out[210]), .A(data_out[202]), .S(shift_en), .Y(n1619)
         );
  INVX1 U1695 ( .A(n1620), .Y(n851) );
  MUX2X1 U1696 ( .B(data_out[218]), .A(data_out[210]), .S(shift_en), .Y(n1620)
         );
  INVX1 U1697 ( .A(n1621), .Y(n849) );
  MUX2X1 U1698 ( .B(data_out[226]), .A(data_out[218]), .S(shift_en), .Y(n1621)
         );
  INVX1 U1699 ( .A(n1622), .Y(n847) );
  MUX2X1 U1700 ( .B(data_out[234]), .A(data_out[226]), .S(shift_en), .Y(n1622)
         );
  INVX1 U1701 ( .A(n1623), .Y(n845) );
  MUX2X1 U1702 ( .B(data_out[242]), .A(data_out[234]), .S(shift_en), .Y(n1623)
         );
  INVX1 U1703 ( .A(n1624), .Y(n843) );
  MUX2X1 U1704 ( .B(data_out[250]), .A(data_out[242]), .S(shift_en), .Y(n1624)
         );
  INVX1 U1705 ( .A(n1625), .Y(n841) );
  MUX2X1 U1706 ( .B(data_out[258]), .A(data_out[250]), .S(shift_en), .Y(n1625)
         );
  INVX1 U1707 ( .A(n1626), .Y(n839) );
  MUX2X1 U1708 ( .B(data_out[266]), .A(data_out[258]), .S(shift_en), .Y(n1626)
         );
  INVX1 U1709 ( .A(n1627), .Y(n837) );
  MUX2X1 U1710 ( .B(data_out[274]), .A(data_out[266]), .S(shift_en), .Y(n1627)
         );
  INVX1 U1711 ( .A(n1628), .Y(n835) );
  MUX2X1 U1712 ( .B(data_out[282]), .A(data_out[274]), .S(shift_en), .Y(n1628)
         );
  INVX1 U1713 ( .A(n1629), .Y(n833) );
  MUX2X1 U1714 ( .B(data_out[290]), .A(data_out[282]), .S(shift_en), .Y(n1629)
         );
  INVX1 U1715 ( .A(n1630), .Y(n831) );
  MUX2X1 U1716 ( .B(data_out[298]), .A(data_out[290]), .S(shift_en), .Y(n1630)
         );
  INVX1 U1717 ( .A(n1631), .Y(n829) );
  MUX2X1 U1718 ( .B(data_out[306]), .A(data_out[298]), .S(shift_en), .Y(n1631)
         );
  INVX1 U1719 ( .A(n1632), .Y(n827) );
  MUX2X1 U1720 ( .B(data_out[314]), .A(data_out[306]), .S(shift_en), .Y(n1632)
         );
  INVX1 U1721 ( .A(n1633), .Y(n825) );
  MUX2X1 U1722 ( .B(data_out[322]), .A(data_out[314]), .S(shift_en), .Y(n1633)
         );
  INVX1 U1723 ( .A(n1634), .Y(n823) );
  MUX2X1 U1724 ( .B(data_out[330]), .A(data_out[322]), .S(shift_en), .Y(n1634)
         );
  INVX1 U1725 ( .A(n1635), .Y(n821) );
  MUX2X1 U1726 ( .B(data_out[338]), .A(data_out[330]), .S(shift_en), .Y(n1635)
         );
  INVX1 U1727 ( .A(n1636), .Y(n819) );
  MUX2X1 U1728 ( .B(data_out[346]), .A(data_out[338]), .S(shift_en), .Y(n1636)
         );
  INVX1 U1729 ( .A(n1637), .Y(n817) );
  MUX2X1 U1730 ( .B(data_out[354]), .A(data_out[346]), .S(shift_en), .Y(n1637)
         );
  INVX1 U1731 ( .A(n1638), .Y(n815) );
  MUX2X1 U1732 ( .B(data_out[362]), .A(data_out[354]), .S(shift_en), .Y(n1638)
         );
  INVX1 U1733 ( .A(n1639), .Y(n813) );
  MUX2X1 U1734 ( .B(data_out[370]), .A(data_out[362]), .S(shift_en), .Y(n1639)
         );
  INVX1 U1735 ( .A(n1640), .Y(n811) );
  MUX2X1 U1736 ( .B(data_out[378]), .A(data_out[370]), .S(shift_en), .Y(n1640)
         );
  INVX1 U1737 ( .A(n1641), .Y(n809) );
  MUX2X1 U1738 ( .B(data_out[386]), .A(data_out[378]), .S(shift_en), .Y(n1641)
         );
  INVX1 U1739 ( .A(n1642), .Y(n807) );
  MUX2X1 U1740 ( .B(data_out[394]), .A(data_out[386]), .S(shift_en), .Y(n1642)
         );
  INVX1 U1741 ( .A(n1643), .Y(n805) );
  MUX2X1 U1742 ( .B(data_out[402]), .A(data_out[394]), .S(shift_en), .Y(n1643)
         );
  INVX1 U1743 ( .A(n1644), .Y(n803) );
  MUX2X1 U1744 ( .B(data_out[410]), .A(data_out[402]), .S(shift_en), .Y(n1644)
         );
  INVX1 U1745 ( .A(n1645), .Y(n801) );
  MUX2X1 U1746 ( .B(data_out[418]), .A(data_out[410]), .S(shift_en), .Y(n1645)
         );
  INVX1 U1747 ( .A(n1646), .Y(n799) );
  MUX2X1 U1748 ( .B(data_out[426]), .A(data_out[418]), .S(shift_en), .Y(n1646)
         );
  INVX1 U1749 ( .A(n1647), .Y(n797) );
  MUX2X1 U1750 ( .B(data_out[434]), .A(data_out[426]), .S(shift_en), .Y(n1647)
         );
  INVX1 U1751 ( .A(n1648), .Y(n795) );
  MUX2X1 U1752 ( .B(data_out[442]), .A(data_out[434]), .S(shift_en), .Y(n1648)
         );
  INVX1 U1753 ( .A(n1649), .Y(n793) );
  MUX2X1 U1754 ( .B(data_out[450]), .A(data_out[442]), .S(shift_en), .Y(n1649)
         );
  INVX1 U1755 ( .A(n1650), .Y(n791) );
  MUX2X1 U1756 ( .B(data_out[458]), .A(data_out[450]), .S(shift_en), .Y(n1650)
         );
  INVX1 U1757 ( .A(n1651), .Y(n789) );
  MUX2X1 U1758 ( .B(data_out[466]), .A(data_out[458]), .S(shift_en), .Y(n1651)
         );
  INVX1 U1759 ( .A(n1652), .Y(n787) );
  MUX2X1 U1760 ( .B(data_out[474]), .A(data_out[466]), .S(shift_en), .Y(n1652)
         );
  INVX1 U1761 ( .A(n1653), .Y(n785) );
  MUX2X1 U1762 ( .B(data_out[482]), .A(data_out[474]), .S(shift_en), .Y(n1653)
         );
  INVX1 U1763 ( .A(n1654), .Y(n783) );
  MUX2X1 U1764 ( .B(data_out[490]), .A(data_out[482]), .S(shift_en), .Y(n1654)
         );
  INVX1 U1765 ( .A(n1655), .Y(n781) );
  MUX2X1 U1766 ( .B(data_out[498]), .A(data_out[490]), .S(shift_en), .Y(n1655)
         );
  INVX1 U1767 ( .A(n1656), .Y(n779) );
  MUX2X1 U1768 ( .B(data_out[506]), .A(data_out[498]), .S(shift_en), .Y(n1656)
         );
  INVX1 U1769 ( .A(n1657), .Y(n777) );
  MUX2X1 U1770 ( .B(data_out[1]), .A(data_in[1]), .S(shift_en), .Y(n1657) );
  INVX1 U1771 ( .A(n1658), .Y(n775) );
  MUX2X1 U1772 ( .B(data_out[9]), .A(data_out[1]), .S(shift_en), .Y(n1658) );
  INVX1 U1773 ( .A(n1659), .Y(n773) );
  MUX2X1 U1774 ( .B(data_out[17]), .A(data_out[9]), .S(shift_en), .Y(n1659) );
  INVX1 U1775 ( .A(n1660), .Y(n771) );
  MUX2X1 U1776 ( .B(data_out[25]), .A(data_out[17]), .S(shift_en), .Y(n1660)
         );
  INVX1 U1777 ( .A(n1661), .Y(n769) );
  MUX2X1 U1778 ( .B(data_out[33]), .A(data_out[25]), .S(shift_en), .Y(n1661)
         );
  INVX1 U1779 ( .A(n1662), .Y(n767) );
  MUX2X1 U1780 ( .B(data_out[41]), .A(data_out[33]), .S(shift_en), .Y(n1662)
         );
  INVX1 U1781 ( .A(n1663), .Y(n765) );
  MUX2X1 U1782 ( .B(data_out[49]), .A(data_out[41]), .S(shift_en), .Y(n1663)
         );
  INVX1 U1783 ( .A(n1664), .Y(n763) );
  MUX2X1 U1784 ( .B(data_out[57]), .A(data_out[49]), .S(shift_en), .Y(n1664)
         );
  INVX1 U1785 ( .A(n1665), .Y(n761) );
  MUX2X1 U1786 ( .B(data_out[65]), .A(data_out[57]), .S(shift_en), .Y(n1665)
         );
  INVX1 U1787 ( .A(n1666), .Y(n759) );
  MUX2X1 U1788 ( .B(data_out[73]), .A(data_out[65]), .S(shift_en), .Y(n1666)
         );
  INVX1 U1789 ( .A(n1667), .Y(n757) );
  MUX2X1 U1790 ( .B(data_out[81]), .A(data_out[73]), .S(shift_en), .Y(n1667)
         );
  INVX1 U1791 ( .A(n1668), .Y(n755) );
  MUX2X1 U1792 ( .B(data_out[89]), .A(data_out[81]), .S(shift_en), .Y(n1668)
         );
  INVX1 U1793 ( .A(n1669), .Y(n753) );
  MUX2X1 U1794 ( .B(data_out[97]), .A(data_out[89]), .S(shift_en), .Y(n1669)
         );
  INVX1 U1795 ( .A(n1670), .Y(n751) );
  MUX2X1 U1796 ( .B(data_out[105]), .A(data_out[97]), .S(shift_en), .Y(n1670)
         );
  INVX1 U1797 ( .A(n1671), .Y(n749) );
  MUX2X1 U1798 ( .B(data_out[113]), .A(data_out[105]), .S(shift_en), .Y(n1671)
         );
  INVX1 U1799 ( .A(n1672), .Y(n747) );
  MUX2X1 U1800 ( .B(data_out[121]), .A(data_out[113]), .S(shift_en), .Y(n1672)
         );
  INVX1 U1801 ( .A(n1673), .Y(n745) );
  MUX2X1 U1802 ( .B(data_out[129]), .A(data_out[121]), .S(shift_en), .Y(n1673)
         );
  INVX1 U1803 ( .A(n1674), .Y(n743) );
  MUX2X1 U1804 ( .B(data_out[137]), .A(data_out[129]), .S(shift_en), .Y(n1674)
         );
  INVX1 U1805 ( .A(n1675), .Y(n741) );
  MUX2X1 U1806 ( .B(data_out[145]), .A(data_out[137]), .S(shift_en), .Y(n1675)
         );
  INVX1 U1807 ( .A(n1676), .Y(n739) );
  MUX2X1 U1808 ( .B(data_out[153]), .A(data_out[145]), .S(shift_en), .Y(n1676)
         );
  INVX1 U1809 ( .A(n1677), .Y(n737) );
  MUX2X1 U1810 ( .B(data_out[161]), .A(data_out[153]), .S(shift_en), .Y(n1677)
         );
  INVX1 U1811 ( .A(n1678), .Y(n735) );
  MUX2X1 U1812 ( .B(data_out[169]), .A(data_out[161]), .S(shift_en), .Y(n1678)
         );
  INVX1 U1813 ( .A(n1679), .Y(n733) );
  MUX2X1 U1814 ( .B(data_out[177]), .A(data_out[169]), .S(shift_en), .Y(n1679)
         );
  INVX1 U1815 ( .A(n1680), .Y(n731) );
  MUX2X1 U1816 ( .B(data_out[185]), .A(data_out[177]), .S(shift_en), .Y(n1680)
         );
  INVX1 U1817 ( .A(n1681), .Y(n729) );
  MUX2X1 U1818 ( .B(data_out[193]), .A(data_out[185]), .S(shift_en), .Y(n1681)
         );
  INVX1 U1819 ( .A(n1682), .Y(n727) );
  MUX2X1 U1820 ( .B(data_out[201]), .A(data_out[193]), .S(shift_en), .Y(n1682)
         );
  INVX1 U1821 ( .A(n1683), .Y(n725) );
  MUX2X1 U1822 ( .B(data_out[209]), .A(data_out[201]), .S(shift_en), .Y(n1683)
         );
  INVX1 U1823 ( .A(n1684), .Y(n723) );
  MUX2X1 U1824 ( .B(data_out[217]), .A(data_out[209]), .S(shift_en), .Y(n1684)
         );
  INVX1 U1825 ( .A(n1685), .Y(n721) );
  MUX2X1 U1826 ( .B(data_out[225]), .A(data_out[217]), .S(shift_en), .Y(n1685)
         );
  INVX1 U1827 ( .A(n1686), .Y(n719) );
  MUX2X1 U1828 ( .B(data_out[233]), .A(data_out[225]), .S(shift_en), .Y(n1686)
         );
  INVX1 U1829 ( .A(n1687), .Y(n717) );
  MUX2X1 U1830 ( .B(data_out[241]), .A(data_out[233]), .S(shift_en), .Y(n1687)
         );
  INVX1 U1831 ( .A(n1688), .Y(n715) );
  MUX2X1 U1832 ( .B(data_out[249]), .A(data_out[241]), .S(shift_en), .Y(n1688)
         );
  INVX1 U1833 ( .A(n1689), .Y(n713) );
  MUX2X1 U1834 ( .B(data_out[257]), .A(data_out[249]), .S(shift_en), .Y(n1689)
         );
  INVX1 U1835 ( .A(n1690), .Y(n711) );
  MUX2X1 U1836 ( .B(data_out[265]), .A(data_out[257]), .S(shift_en), .Y(n1690)
         );
  INVX1 U1837 ( .A(n1691), .Y(n709) );
  MUX2X1 U1838 ( .B(data_out[273]), .A(data_out[265]), .S(shift_en), .Y(n1691)
         );
  INVX1 U1839 ( .A(n1692), .Y(n707) );
  MUX2X1 U1840 ( .B(data_out[281]), .A(data_out[273]), .S(shift_en), .Y(n1692)
         );
  INVX1 U1841 ( .A(n1693), .Y(n705) );
  MUX2X1 U1842 ( .B(data_out[289]), .A(data_out[281]), .S(shift_en), .Y(n1693)
         );
  INVX1 U1843 ( .A(n1694), .Y(n703) );
  MUX2X1 U1844 ( .B(data_out[297]), .A(data_out[289]), .S(shift_en), .Y(n1694)
         );
  INVX1 U1845 ( .A(n1695), .Y(n701) );
  MUX2X1 U1846 ( .B(data_out[305]), .A(data_out[297]), .S(shift_en), .Y(n1695)
         );
  INVX1 U1847 ( .A(n1696), .Y(n699) );
  MUX2X1 U1848 ( .B(data_out[313]), .A(data_out[305]), .S(shift_en), .Y(n1696)
         );
  INVX1 U1849 ( .A(n1697), .Y(n697) );
  MUX2X1 U1850 ( .B(data_out[321]), .A(data_out[313]), .S(shift_en), .Y(n1697)
         );
  INVX1 U1851 ( .A(n1698), .Y(n695) );
  MUX2X1 U1852 ( .B(data_out[329]), .A(data_out[321]), .S(shift_en), .Y(n1698)
         );
  INVX1 U1853 ( .A(n1699), .Y(n693) );
  MUX2X1 U1854 ( .B(data_out[337]), .A(data_out[329]), .S(shift_en), .Y(n1699)
         );
  INVX1 U1855 ( .A(n1700), .Y(n691) );
  MUX2X1 U1856 ( .B(data_out[345]), .A(data_out[337]), .S(shift_en), .Y(n1700)
         );
  INVX1 U1857 ( .A(n1701), .Y(n689) );
  MUX2X1 U1858 ( .B(data_out[353]), .A(data_out[345]), .S(shift_en), .Y(n1701)
         );
  INVX1 U1859 ( .A(n1702), .Y(n687) );
  MUX2X1 U1860 ( .B(data_out[361]), .A(data_out[353]), .S(shift_en), .Y(n1702)
         );
  INVX1 U1861 ( .A(n1703), .Y(n685) );
  MUX2X1 U1862 ( .B(data_out[369]), .A(data_out[361]), .S(shift_en), .Y(n1703)
         );
  INVX1 U1863 ( .A(n1704), .Y(n683) );
  MUX2X1 U1864 ( .B(data_out[377]), .A(data_out[369]), .S(shift_en), .Y(n1704)
         );
  INVX1 U1865 ( .A(n1705), .Y(n681) );
  MUX2X1 U1866 ( .B(data_out[385]), .A(data_out[377]), .S(shift_en), .Y(n1705)
         );
  INVX1 U1867 ( .A(n1706), .Y(n679) );
  MUX2X1 U1868 ( .B(data_out[393]), .A(data_out[385]), .S(shift_en), .Y(n1706)
         );
  INVX1 U1869 ( .A(n1707), .Y(n677) );
  MUX2X1 U1870 ( .B(data_out[401]), .A(data_out[393]), .S(shift_en), .Y(n1707)
         );
  INVX1 U1871 ( .A(n1708), .Y(n675) );
  MUX2X1 U1872 ( .B(data_out[409]), .A(data_out[401]), .S(shift_en), .Y(n1708)
         );
  INVX1 U1873 ( .A(n1709), .Y(n673) );
  MUX2X1 U1874 ( .B(data_out[417]), .A(data_out[409]), .S(shift_en), .Y(n1709)
         );
  INVX1 U1875 ( .A(n1710), .Y(n671) );
  MUX2X1 U1876 ( .B(data_out[425]), .A(data_out[417]), .S(shift_en), .Y(n1710)
         );
  INVX1 U1877 ( .A(n1711), .Y(n669) );
  MUX2X1 U1878 ( .B(data_out[433]), .A(data_out[425]), .S(shift_en), .Y(n1711)
         );
  INVX1 U1879 ( .A(n1712), .Y(n667) );
  MUX2X1 U1880 ( .B(data_out[441]), .A(data_out[433]), .S(shift_en), .Y(n1712)
         );
  INVX1 U1881 ( .A(n1713), .Y(n665) );
  MUX2X1 U1882 ( .B(data_out[449]), .A(data_out[441]), .S(shift_en), .Y(n1713)
         );
  INVX1 U1883 ( .A(n1714), .Y(n663) );
  MUX2X1 U1884 ( .B(data_out[457]), .A(data_out[449]), .S(shift_en), .Y(n1714)
         );
  INVX1 U1885 ( .A(n1715), .Y(n661) );
  MUX2X1 U1886 ( .B(data_out[465]), .A(data_out[457]), .S(shift_en), .Y(n1715)
         );
  INVX1 U1887 ( .A(n1716), .Y(n659) );
  MUX2X1 U1888 ( .B(data_out[473]), .A(data_out[465]), .S(shift_en), .Y(n1716)
         );
  INVX1 U1889 ( .A(n1717), .Y(n657) );
  MUX2X1 U1890 ( .B(data_out[481]), .A(data_out[473]), .S(shift_en), .Y(n1717)
         );
  INVX1 U1891 ( .A(n1718), .Y(n655) );
  MUX2X1 U1892 ( .B(data_out[489]), .A(data_out[481]), .S(shift_en), .Y(n1718)
         );
  INVX1 U1893 ( .A(n1719), .Y(n653) );
  MUX2X1 U1894 ( .B(data_out[497]), .A(data_out[489]), .S(shift_en), .Y(n1719)
         );
  INVX1 U1895 ( .A(n1720), .Y(n651) );
  MUX2X1 U1896 ( .B(data_out[505]), .A(data_out[497]), .S(shift_en), .Y(n1720)
         );
  INVX1 U1897 ( .A(n1721), .Y(n649) );
  MUX2X1 U1898 ( .B(data_out[0]), .A(data_in[0]), .S(shift_en), .Y(n1721) );
  INVX1 U1899 ( .A(n1722), .Y(n647) );
  MUX2X1 U1900 ( .B(data_out[8]), .A(data_out[0]), .S(shift_en), .Y(n1722) );
  INVX1 U1901 ( .A(n1723), .Y(n645) );
  MUX2X1 U1902 ( .B(data_out[16]), .A(data_out[8]), .S(shift_en), .Y(n1723) );
  INVX1 U1903 ( .A(n1724), .Y(n643) );
  MUX2X1 U1904 ( .B(data_out[24]), .A(data_out[16]), .S(shift_en), .Y(n1724)
         );
  INVX1 U1905 ( .A(n1725), .Y(n641) );
  MUX2X1 U1906 ( .B(data_out[32]), .A(data_out[24]), .S(shift_en), .Y(n1725)
         );
  INVX1 U1907 ( .A(n1726), .Y(n639) );
  MUX2X1 U1908 ( .B(data_out[40]), .A(data_out[32]), .S(shift_en), .Y(n1726)
         );
  INVX1 U1909 ( .A(n1727), .Y(n637) );
  MUX2X1 U1910 ( .B(data_out[48]), .A(data_out[40]), .S(shift_en), .Y(n1727)
         );
  INVX1 U1911 ( .A(n1728), .Y(n635) );
  MUX2X1 U1912 ( .B(data_out[56]), .A(data_out[48]), .S(shift_en), .Y(n1728)
         );
  INVX1 U1913 ( .A(n1729), .Y(n633) );
  MUX2X1 U1914 ( .B(data_out[64]), .A(data_out[56]), .S(shift_en), .Y(n1729)
         );
  INVX1 U1915 ( .A(n1730), .Y(n631) );
  MUX2X1 U1916 ( .B(data_out[72]), .A(data_out[64]), .S(shift_en), .Y(n1730)
         );
  INVX1 U1917 ( .A(n1731), .Y(n629) );
  MUX2X1 U1918 ( .B(data_out[80]), .A(data_out[72]), .S(shift_en), .Y(n1731)
         );
  INVX1 U1919 ( .A(n1732), .Y(n627) );
  MUX2X1 U1920 ( .B(data_out[88]), .A(data_out[80]), .S(shift_en), .Y(n1732)
         );
  INVX1 U1921 ( .A(n1733), .Y(n625) );
  MUX2X1 U1922 ( .B(data_out[96]), .A(data_out[88]), .S(shift_en), .Y(n1733)
         );
  INVX1 U1923 ( .A(n1734), .Y(n623) );
  MUX2X1 U1924 ( .B(data_out[104]), .A(data_out[96]), .S(shift_en), .Y(n1734)
         );
  INVX1 U1925 ( .A(n1735), .Y(n621) );
  MUX2X1 U1926 ( .B(data_out[112]), .A(data_out[104]), .S(shift_en), .Y(n1735)
         );
  INVX1 U1927 ( .A(n1736), .Y(n619) );
  MUX2X1 U1928 ( .B(data_out[120]), .A(data_out[112]), .S(shift_en), .Y(n1736)
         );
  INVX1 U1929 ( .A(n1737), .Y(n617) );
  MUX2X1 U1930 ( .B(data_out[128]), .A(data_out[120]), .S(shift_en), .Y(n1737)
         );
  INVX1 U1931 ( .A(n1738), .Y(n615) );
  MUX2X1 U1932 ( .B(data_out[136]), .A(data_out[128]), .S(shift_en), .Y(n1738)
         );
  INVX1 U1933 ( .A(n1739), .Y(n613) );
  MUX2X1 U1934 ( .B(data_out[144]), .A(data_out[136]), .S(shift_en), .Y(n1739)
         );
  INVX1 U1935 ( .A(n1740), .Y(n611) );
  MUX2X1 U1936 ( .B(data_out[152]), .A(data_out[144]), .S(shift_en), .Y(n1740)
         );
  INVX1 U1937 ( .A(n1741), .Y(n609) );
  MUX2X1 U1938 ( .B(data_out[160]), .A(data_out[152]), .S(shift_en), .Y(n1741)
         );
  INVX1 U1939 ( .A(n1742), .Y(n607) );
  MUX2X1 U1940 ( .B(data_out[168]), .A(data_out[160]), .S(shift_en), .Y(n1742)
         );
  INVX1 U1941 ( .A(n1743), .Y(n605) );
  MUX2X1 U1942 ( .B(data_out[176]), .A(data_out[168]), .S(shift_en), .Y(n1743)
         );
  INVX1 U1943 ( .A(n1744), .Y(n603) );
  MUX2X1 U1944 ( .B(data_out[184]), .A(data_out[176]), .S(shift_en), .Y(n1744)
         );
  INVX1 U1945 ( .A(n1745), .Y(n601) );
  MUX2X1 U1946 ( .B(data_out[192]), .A(data_out[184]), .S(shift_en), .Y(n1745)
         );
  INVX1 U1947 ( .A(n1746), .Y(n599) );
  MUX2X1 U1948 ( .B(data_out[200]), .A(data_out[192]), .S(shift_en), .Y(n1746)
         );
  INVX1 U1949 ( .A(n1747), .Y(n597) );
  MUX2X1 U1950 ( .B(data_out[208]), .A(data_out[200]), .S(shift_en), .Y(n1747)
         );
  INVX1 U1951 ( .A(n1748), .Y(n595) );
  MUX2X1 U1952 ( .B(data_out[216]), .A(data_out[208]), .S(shift_en), .Y(n1748)
         );
  INVX1 U1953 ( .A(n1749), .Y(n593) );
  MUX2X1 U1954 ( .B(data_out[224]), .A(data_out[216]), .S(shift_en), .Y(n1749)
         );
  INVX1 U1955 ( .A(n1750), .Y(n591) );
  MUX2X1 U1956 ( .B(data_out[232]), .A(data_out[224]), .S(shift_en), .Y(n1750)
         );
  INVX1 U1957 ( .A(n1751), .Y(n589) );
  MUX2X1 U1958 ( .B(data_out[240]), .A(data_out[232]), .S(shift_en), .Y(n1751)
         );
  INVX1 U1959 ( .A(n1752), .Y(n587) );
  MUX2X1 U1960 ( .B(data_out[248]), .A(data_out[240]), .S(shift_en), .Y(n1752)
         );
  INVX1 U1961 ( .A(n1753), .Y(n585) );
  MUX2X1 U1962 ( .B(data_out[256]), .A(data_out[248]), .S(shift_en), .Y(n1753)
         );
  INVX1 U1963 ( .A(n1754), .Y(n583) );
  MUX2X1 U1964 ( .B(data_out[264]), .A(data_out[256]), .S(shift_en), .Y(n1754)
         );
  INVX1 U1965 ( .A(n1755), .Y(n581) );
  MUX2X1 U1966 ( .B(data_out[272]), .A(data_out[264]), .S(shift_en), .Y(n1755)
         );
  INVX1 U1967 ( .A(n1756), .Y(n579) );
  MUX2X1 U1968 ( .B(data_out[280]), .A(data_out[272]), .S(shift_en), .Y(n1756)
         );
  INVX1 U1969 ( .A(n1757), .Y(n577) );
  MUX2X1 U1970 ( .B(data_out[288]), .A(data_out[280]), .S(shift_en), .Y(n1757)
         );
  INVX1 U1971 ( .A(n1758), .Y(n575) );
  MUX2X1 U1972 ( .B(data_out[296]), .A(data_out[288]), .S(shift_en), .Y(n1758)
         );
  INVX1 U1973 ( .A(n1759), .Y(n573) );
  MUX2X1 U1974 ( .B(data_out[304]), .A(data_out[296]), .S(shift_en), .Y(n1759)
         );
  INVX1 U1975 ( .A(n1760), .Y(n571) );
  MUX2X1 U1976 ( .B(data_out[312]), .A(data_out[304]), .S(shift_en), .Y(n1760)
         );
  INVX1 U1977 ( .A(n1761), .Y(n569) );
  MUX2X1 U1978 ( .B(data_out[320]), .A(data_out[312]), .S(shift_en), .Y(n1761)
         );
  INVX1 U1979 ( .A(n1762), .Y(n567) );
  MUX2X1 U1980 ( .B(data_out[328]), .A(data_out[320]), .S(shift_en), .Y(n1762)
         );
  INVX1 U1981 ( .A(n1763), .Y(n565) );
  MUX2X1 U1982 ( .B(data_out[336]), .A(data_out[328]), .S(shift_en), .Y(n1763)
         );
  INVX1 U1983 ( .A(n1764), .Y(n563) );
  MUX2X1 U1984 ( .B(data_out[344]), .A(data_out[336]), .S(shift_en), .Y(n1764)
         );
  INVX1 U1985 ( .A(n1765), .Y(n561) );
  MUX2X1 U1986 ( .B(data_out[352]), .A(data_out[344]), .S(shift_en), .Y(n1765)
         );
  INVX1 U1987 ( .A(n1766), .Y(n559) );
  MUX2X1 U1988 ( .B(data_out[360]), .A(data_out[352]), .S(shift_en), .Y(n1766)
         );
  INVX1 U1989 ( .A(n1767), .Y(n557) );
  MUX2X1 U1990 ( .B(data_out[368]), .A(data_out[360]), .S(shift_en), .Y(n1767)
         );
  INVX1 U1991 ( .A(n1768), .Y(n555) );
  MUX2X1 U1992 ( .B(data_out[376]), .A(data_out[368]), .S(shift_en), .Y(n1768)
         );
  INVX1 U1993 ( .A(n1769), .Y(n553) );
  MUX2X1 U1994 ( .B(data_out[384]), .A(data_out[376]), .S(shift_en), .Y(n1769)
         );
  INVX1 U1995 ( .A(n1770), .Y(n551) );
  MUX2X1 U1996 ( .B(data_out[392]), .A(data_out[384]), .S(shift_en), .Y(n1770)
         );
  INVX1 U1997 ( .A(n1771), .Y(n549) );
  MUX2X1 U1998 ( .B(data_out[400]), .A(data_out[392]), .S(shift_en), .Y(n1771)
         );
  INVX1 U1999 ( .A(n1772), .Y(n547) );
  MUX2X1 U2000 ( .B(data_out[408]), .A(data_out[400]), .S(shift_en), .Y(n1772)
         );
  INVX1 U2001 ( .A(n1773), .Y(n545) );
  MUX2X1 U2002 ( .B(data_out[416]), .A(data_out[408]), .S(shift_en), .Y(n1773)
         );
  INVX1 U2003 ( .A(n1774), .Y(n543) );
  MUX2X1 U2004 ( .B(data_out[424]), .A(data_out[416]), .S(shift_en), .Y(n1774)
         );
  INVX1 U2005 ( .A(n1775), .Y(n541) );
  MUX2X1 U2006 ( .B(data_out[432]), .A(data_out[424]), .S(shift_en), .Y(n1775)
         );
  INVX1 U2007 ( .A(n1776), .Y(n539) );
  MUX2X1 U2008 ( .B(data_out[440]), .A(data_out[432]), .S(shift_en), .Y(n1776)
         );
  INVX1 U2009 ( .A(n1777), .Y(n537) );
  MUX2X1 U2010 ( .B(data_out[448]), .A(data_out[440]), .S(shift_en), .Y(n1777)
         );
  INVX1 U2011 ( .A(n1778), .Y(n535) );
  MUX2X1 U2012 ( .B(data_out[456]), .A(data_out[448]), .S(shift_en), .Y(n1778)
         );
  INVX1 U2013 ( .A(n1779), .Y(n533) );
  MUX2X1 U2014 ( .B(data_out[464]), .A(data_out[456]), .S(shift_en), .Y(n1779)
         );
  INVX1 U2015 ( .A(n1780), .Y(n531) );
  MUX2X1 U2016 ( .B(data_out[472]), .A(data_out[464]), .S(shift_en), .Y(n1780)
         );
  INVX1 U2017 ( .A(n1781), .Y(n529) );
  MUX2X1 U2018 ( .B(data_out[480]), .A(data_out[472]), .S(shift_en), .Y(n1781)
         );
  INVX1 U2019 ( .A(n1782), .Y(n527) );
  MUX2X1 U2020 ( .B(data_out[488]), .A(data_out[480]), .S(shift_en), .Y(n1782)
         );
  INVX1 U2021 ( .A(n1783), .Y(n525) );
  MUX2X1 U2022 ( .B(data_out[496]), .A(data_out[488]), .S(shift_en), .Y(n1783)
         );
  INVX1 U2023 ( .A(n1784), .Y(n523) );
  MUX2X1 U2024 ( .B(data_out[504]), .A(data_out[496]), .S(shift_en), .Y(n1784)
         );
  INVX1 U2025 ( .A(n1785), .Y(n1545) );
  MUX2X1 U2026 ( .B(data_out[7]), .A(data_in[7]), .S(shift_en), .Y(n1785) );
  INVX1 U2027 ( .A(n1786), .Y(n1543) );
  MUX2X1 U2028 ( .B(data_out[15]), .A(data_out[7]), .S(shift_en), .Y(n1786) );
  INVX1 U2029 ( .A(n1787), .Y(n1541) );
  MUX2X1 U2030 ( .B(data_out[23]), .A(data_out[15]), .S(shift_en), .Y(n1787)
         );
  INVX1 U2031 ( .A(n1788), .Y(n1539) );
  MUX2X1 U2032 ( .B(data_out[31]), .A(data_out[23]), .S(shift_en), .Y(n1788)
         );
  INVX1 U2033 ( .A(n1789), .Y(n1537) );
  MUX2X1 U2034 ( .B(data_out[39]), .A(data_out[31]), .S(shift_en), .Y(n1789)
         );
  INVX1 U2035 ( .A(n1790), .Y(n1535) );
  MUX2X1 U2036 ( .B(data_out[47]), .A(data_out[39]), .S(shift_en), .Y(n1790)
         );
  INVX1 U2037 ( .A(n1791), .Y(n1533) );
  MUX2X1 U2038 ( .B(data_out[55]), .A(data_out[47]), .S(shift_en), .Y(n1791)
         );
  INVX1 U2039 ( .A(n1792), .Y(n1531) );
  MUX2X1 U2040 ( .B(data_out[63]), .A(data_out[55]), .S(shift_en), .Y(n1792)
         );
  INVX1 U2041 ( .A(n1793), .Y(n1529) );
  MUX2X1 U2042 ( .B(data_out[71]), .A(data_out[63]), .S(shift_en), .Y(n1793)
         );
  INVX1 U2043 ( .A(n1794), .Y(n1527) );
  MUX2X1 U2044 ( .B(data_out[79]), .A(data_out[71]), .S(shift_en), .Y(n1794)
         );
  INVX1 U2045 ( .A(n1795), .Y(n1525) );
  MUX2X1 U2046 ( .B(data_out[87]), .A(data_out[79]), .S(shift_en), .Y(n1795)
         );
  INVX1 U2047 ( .A(n1796), .Y(n1523) );
  MUX2X1 U2048 ( .B(data_out[95]), .A(data_out[87]), .S(shift_en), .Y(n1796)
         );
  INVX1 U2049 ( .A(n1797), .Y(n1521) );
  MUX2X1 U2050 ( .B(data_out[103]), .A(data_out[95]), .S(shift_en), .Y(n1797)
         );
  INVX1 U2051 ( .A(n1798), .Y(n1519) );
  MUX2X1 U2052 ( .B(data_out[111]), .A(data_out[103]), .S(shift_en), .Y(n1798)
         );
  INVX1 U2053 ( .A(n1799), .Y(n1517) );
  MUX2X1 U2054 ( .B(data_out[119]), .A(data_out[111]), .S(shift_en), .Y(n1799)
         );
  INVX1 U2055 ( .A(n1800), .Y(n1515) );
  MUX2X1 U2056 ( .B(data_out[127]), .A(data_out[119]), .S(shift_en), .Y(n1800)
         );
  INVX1 U2057 ( .A(n1801), .Y(n1513) );
  MUX2X1 U2058 ( .B(data_out[135]), .A(data_out[127]), .S(shift_en), .Y(n1801)
         );
  INVX1 U2059 ( .A(n1802), .Y(n1511) );
  MUX2X1 U2060 ( .B(data_out[143]), .A(data_out[135]), .S(shift_en), .Y(n1802)
         );
  INVX1 U2061 ( .A(n1803), .Y(n1509) );
  MUX2X1 U2062 ( .B(data_out[151]), .A(data_out[143]), .S(shift_en), .Y(n1803)
         );
  INVX1 U2063 ( .A(n1804), .Y(n1507) );
  MUX2X1 U2064 ( .B(data_out[159]), .A(data_out[151]), .S(shift_en), .Y(n1804)
         );
  INVX1 U2065 ( .A(n1805), .Y(n1505) );
  MUX2X1 U2066 ( .B(data_out[167]), .A(data_out[159]), .S(shift_en), .Y(n1805)
         );
  INVX1 U2067 ( .A(n1806), .Y(n1503) );
  MUX2X1 U2068 ( .B(data_out[175]), .A(data_out[167]), .S(shift_en), .Y(n1806)
         );
  INVX1 U2069 ( .A(n1807), .Y(n1501) );
  MUX2X1 U2070 ( .B(data_out[183]), .A(data_out[175]), .S(shift_en), .Y(n1807)
         );
  INVX1 U2071 ( .A(n1808), .Y(n1499) );
  MUX2X1 U2072 ( .B(data_out[191]), .A(data_out[183]), .S(shift_en), .Y(n1808)
         );
  INVX1 U2073 ( .A(n1809), .Y(n1497) );
  MUX2X1 U2074 ( .B(data_out[199]), .A(data_out[191]), .S(shift_en), .Y(n1809)
         );
  INVX1 U2075 ( .A(n1810), .Y(n1495) );
  MUX2X1 U2076 ( .B(data_out[207]), .A(data_out[199]), .S(shift_en), .Y(n1810)
         );
  INVX1 U2077 ( .A(n1811), .Y(n1493) );
  MUX2X1 U2078 ( .B(data_out[215]), .A(data_out[207]), .S(shift_en), .Y(n1811)
         );
  INVX1 U2079 ( .A(n1812), .Y(n1491) );
  MUX2X1 U2080 ( .B(data_out[223]), .A(data_out[215]), .S(shift_en), .Y(n1812)
         );
  INVX1 U2081 ( .A(n1813), .Y(n1489) );
  MUX2X1 U2082 ( .B(data_out[231]), .A(data_out[223]), .S(shift_en), .Y(n1813)
         );
  INVX1 U2083 ( .A(n1814), .Y(n1487) );
  MUX2X1 U2084 ( .B(data_out[239]), .A(data_out[231]), .S(shift_en), .Y(n1814)
         );
  INVX1 U2085 ( .A(n1815), .Y(n1485) );
  MUX2X1 U2086 ( .B(data_out[247]), .A(data_out[239]), .S(shift_en), .Y(n1815)
         );
  INVX1 U2087 ( .A(n1816), .Y(n1483) );
  MUX2X1 U2088 ( .B(data_out[255]), .A(data_out[247]), .S(shift_en), .Y(n1816)
         );
  INVX1 U2089 ( .A(n1817), .Y(n1481) );
  MUX2X1 U2090 ( .B(data_out[263]), .A(data_out[255]), .S(shift_en), .Y(n1817)
         );
  INVX1 U2091 ( .A(n1818), .Y(n1479) );
  MUX2X1 U2092 ( .B(data_out[271]), .A(data_out[263]), .S(shift_en), .Y(n1818)
         );
  INVX1 U2093 ( .A(n1819), .Y(n1477) );
  MUX2X1 U2094 ( .B(data_out[279]), .A(data_out[271]), .S(shift_en), .Y(n1819)
         );
  INVX1 U2095 ( .A(n1820), .Y(n1475) );
  MUX2X1 U2096 ( .B(data_out[287]), .A(data_out[279]), .S(shift_en), .Y(n1820)
         );
  INVX1 U2097 ( .A(n1821), .Y(n1473) );
  MUX2X1 U2098 ( .B(data_out[295]), .A(data_out[287]), .S(shift_en), .Y(n1821)
         );
  INVX1 U2099 ( .A(n1822), .Y(n1471) );
  MUX2X1 U2100 ( .B(data_out[303]), .A(data_out[295]), .S(shift_en), .Y(n1822)
         );
  INVX1 U2101 ( .A(n1823), .Y(n1469) );
  MUX2X1 U2102 ( .B(data_out[311]), .A(data_out[303]), .S(shift_en), .Y(n1823)
         );
  INVX1 U2103 ( .A(n1824), .Y(n1467) );
  MUX2X1 U2104 ( .B(data_out[319]), .A(data_out[311]), .S(shift_en), .Y(n1824)
         );
  INVX1 U2105 ( .A(n1825), .Y(n1465) );
  MUX2X1 U2106 ( .B(data_out[327]), .A(data_out[319]), .S(shift_en), .Y(n1825)
         );
  INVX1 U2107 ( .A(n1826), .Y(n1463) );
  MUX2X1 U2108 ( .B(data_out[335]), .A(data_out[327]), .S(shift_en), .Y(n1826)
         );
  INVX1 U2109 ( .A(n1827), .Y(n1461) );
  MUX2X1 U2110 ( .B(data_out[343]), .A(data_out[335]), .S(shift_en), .Y(n1827)
         );
  INVX1 U2111 ( .A(n1828), .Y(n1459) );
  MUX2X1 U2112 ( .B(data_out[351]), .A(data_out[343]), .S(shift_en), .Y(n1828)
         );
  INVX1 U2113 ( .A(n1829), .Y(n1457) );
  MUX2X1 U2114 ( .B(data_out[359]), .A(data_out[351]), .S(shift_en), .Y(n1829)
         );
  INVX1 U2115 ( .A(n1830), .Y(n1455) );
  MUX2X1 U2116 ( .B(data_out[367]), .A(data_out[359]), .S(shift_en), .Y(n1830)
         );
  INVX1 U2117 ( .A(n1831), .Y(n1453) );
  MUX2X1 U2118 ( .B(data_out[375]), .A(data_out[367]), .S(shift_en), .Y(n1831)
         );
  INVX1 U2119 ( .A(n1832), .Y(n1451) );
  MUX2X1 U2120 ( .B(data_out[383]), .A(data_out[375]), .S(shift_en), .Y(n1832)
         );
  INVX1 U2121 ( .A(n1833), .Y(n1449) );
  MUX2X1 U2122 ( .B(data_out[391]), .A(data_out[383]), .S(shift_en), .Y(n1833)
         );
  INVX1 U2123 ( .A(n1834), .Y(n1447) );
  MUX2X1 U2124 ( .B(data_out[399]), .A(data_out[391]), .S(shift_en), .Y(n1834)
         );
  INVX1 U2125 ( .A(n1835), .Y(n1445) );
  MUX2X1 U2126 ( .B(data_out[407]), .A(data_out[399]), .S(shift_en), .Y(n1835)
         );
  INVX1 U2127 ( .A(n1836), .Y(n1443) );
  MUX2X1 U2128 ( .B(data_out[415]), .A(data_out[407]), .S(shift_en), .Y(n1836)
         );
  INVX1 U2129 ( .A(n1837), .Y(n1441) );
  MUX2X1 U2130 ( .B(data_out[423]), .A(data_out[415]), .S(shift_en), .Y(n1837)
         );
  INVX1 U2131 ( .A(n1838), .Y(n1439) );
  MUX2X1 U2132 ( .B(data_out[431]), .A(data_out[423]), .S(shift_en), .Y(n1838)
         );
  INVX1 U2133 ( .A(n1839), .Y(n1437) );
  MUX2X1 U2134 ( .B(data_out[439]), .A(data_out[431]), .S(shift_en), .Y(n1839)
         );
  INVX1 U2135 ( .A(n1840), .Y(n1435) );
  MUX2X1 U2136 ( .B(data_out[447]), .A(data_out[439]), .S(shift_en), .Y(n1840)
         );
  INVX1 U2137 ( .A(n1841), .Y(n1433) );
  MUX2X1 U2138 ( .B(data_out[455]), .A(data_out[447]), .S(shift_en), .Y(n1841)
         );
  INVX1 U2139 ( .A(n1842), .Y(n1431) );
  MUX2X1 U2140 ( .B(data_out[463]), .A(data_out[455]), .S(shift_en), .Y(n1842)
         );
  INVX1 U2141 ( .A(n1843), .Y(n1429) );
  MUX2X1 U2142 ( .B(data_out[471]), .A(data_out[463]), .S(shift_en), .Y(n1843)
         );
  INVX1 U2143 ( .A(n1844), .Y(n1427) );
  MUX2X1 U2144 ( .B(data_out[479]), .A(data_out[471]), .S(shift_en), .Y(n1844)
         );
  INVX1 U2145 ( .A(n1845), .Y(n1425) );
  MUX2X1 U2146 ( .B(data_out[487]), .A(data_out[479]), .S(shift_en), .Y(n1845)
         );
  INVX1 U2147 ( .A(n1846), .Y(n1423) );
  MUX2X1 U2148 ( .B(data_out[495]), .A(data_out[487]), .S(shift_en), .Y(n1846)
         );
  INVX1 U2149 ( .A(n1847), .Y(n1421) );
  MUX2X1 U2150 ( .B(data_out[503]), .A(data_out[495]), .S(shift_en), .Y(n1847)
         );
  INVX1 U2151 ( .A(n1848), .Y(n1419) );
  MUX2X1 U2152 ( .B(data_out[511]), .A(data_out[503]), .S(shift_en), .Y(n1848)
         );
  INVX1 U2153 ( .A(n1849), .Y(n1417) );
  MUX2X1 U2154 ( .B(data_out[6]), .A(data_in[6]), .S(shift_en), .Y(n1849) );
  INVX1 U2155 ( .A(n1850), .Y(n1415) );
  MUX2X1 U2156 ( .B(data_out[14]), .A(data_out[6]), .S(shift_en), .Y(n1850) );
  INVX1 U2157 ( .A(n1851), .Y(n1413) );
  MUX2X1 U2158 ( .B(data_out[22]), .A(data_out[14]), .S(shift_en), .Y(n1851)
         );
  INVX1 U2159 ( .A(n1852), .Y(n1411) );
  MUX2X1 U2160 ( .B(data_out[30]), .A(data_out[22]), .S(shift_en), .Y(n1852)
         );
  INVX1 U2161 ( .A(n1853), .Y(n1409) );
  MUX2X1 U2162 ( .B(data_out[38]), .A(data_out[30]), .S(shift_en), .Y(n1853)
         );
  INVX1 U2163 ( .A(n1854), .Y(n1407) );
  MUX2X1 U2164 ( .B(data_out[46]), .A(data_out[38]), .S(shift_en), .Y(n1854)
         );
  INVX1 U2165 ( .A(n1855), .Y(n1405) );
  MUX2X1 U2166 ( .B(data_out[54]), .A(data_out[46]), .S(shift_en), .Y(n1855)
         );
  INVX1 U2167 ( .A(n1856), .Y(n1403) );
  MUX2X1 U2168 ( .B(data_out[62]), .A(data_out[54]), .S(shift_en), .Y(n1856)
         );
  INVX1 U2169 ( .A(n1857), .Y(n1401) );
  MUX2X1 U2170 ( .B(data_out[70]), .A(data_out[62]), .S(shift_en), .Y(n1857)
         );
  INVX1 U2171 ( .A(n1858), .Y(n1399) );
  MUX2X1 U2172 ( .B(data_out[78]), .A(data_out[70]), .S(shift_en), .Y(n1858)
         );
  INVX1 U2173 ( .A(n1859), .Y(n1397) );
  MUX2X1 U2174 ( .B(data_out[86]), .A(data_out[78]), .S(shift_en), .Y(n1859)
         );
  INVX1 U2175 ( .A(n1860), .Y(n1395) );
  MUX2X1 U2176 ( .B(data_out[94]), .A(data_out[86]), .S(shift_en), .Y(n1860)
         );
  INVX1 U2177 ( .A(n1861), .Y(n1393) );
  MUX2X1 U2178 ( .B(data_out[102]), .A(data_out[94]), .S(shift_en), .Y(n1861)
         );
  INVX1 U2179 ( .A(n1862), .Y(n1391) );
  MUX2X1 U2180 ( .B(data_out[110]), .A(data_out[102]), .S(shift_en), .Y(n1862)
         );
  INVX1 U2181 ( .A(n1863), .Y(n1389) );
  MUX2X1 U2182 ( .B(data_out[118]), .A(data_out[110]), .S(shift_en), .Y(n1863)
         );
  INVX1 U2183 ( .A(n1864), .Y(n1387) );
  MUX2X1 U2184 ( .B(data_out[126]), .A(data_out[118]), .S(shift_en), .Y(n1864)
         );
  INVX1 U2185 ( .A(n1865), .Y(n1385) );
  MUX2X1 U2186 ( .B(data_out[134]), .A(data_out[126]), .S(shift_en), .Y(n1865)
         );
  INVX1 U2187 ( .A(n1866), .Y(n1383) );
  MUX2X1 U2188 ( .B(data_out[142]), .A(data_out[134]), .S(shift_en), .Y(n1866)
         );
  INVX1 U2189 ( .A(n1867), .Y(n1381) );
  MUX2X1 U2190 ( .B(data_out[150]), .A(data_out[142]), .S(shift_en), .Y(n1867)
         );
  INVX1 U2191 ( .A(n1868), .Y(n1379) );
  MUX2X1 U2192 ( .B(data_out[158]), .A(data_out[150]), .S(shift_en), .Y(n1868)
         );
  INVX1 U2193 ( .A(n1869), .Y(n1377) );
  MUX2X1 U2194 ( .B(data_out[166]), .A(data_out[158]), .S(shift_en), .Y(n1869)
         );
  INVX1 U2195 ( .A(n1870), .Y(n1375) );
  MUX2X1 U2196 ( .B(data_out[174]), .A(data_out[166]), .S(shift_en), .Y(n1870)
         );
  INVX1 U2197 ( .A(n1871), .Y(n1373) );
  MUX2X1 U2198 ( .B(data_out[182]), .A(data_out[174]), .S(shift_en), .Y(n1871)
         );
  INVX1 U2199 ( .A(n1872), .Y(n1371) );
  MUX2X1 U2200 ( .B(data_out[190]), .A(data_out[182]), .S(shift_en), .Y(n1872)
         );
  INVX1 U2201 ( .A(n1873), .Y(n1369) );
  MUX2X1 U2202 ( .B(data_out[198]), .A(data_out[190]), .S(shift_en), .Y(n1873)
         );
  INVX1 U2203 ( .A(n1874), .Y(n1367) );
  MUX2X1 U2204 ( .B(data_out[206]), .A(data_out[198]), .S(shift_en), .Y(n1874)
         );
  INVX1 U2205 ( .A(n1875), .Y(n1365) );
  MUX2X1 U2206 ( .B(data_out[214]), .A(data_out[206]), .S(shift_en), .Y(n1875)
         );
  INVX1 U2207 ( .A(n1876), .Y(n1363) );
  MUX2X1 U2208 ( .B(data_out[222]), .A(data_out[214]), .S(shift_en), .Y(n1876)
         );
  INVX1 U2209 ( .A(n1877), .Y(n1361) );
  MUX2X1 U2210 ( .B(data_out[230]), .A(data_out[222]), .S(shift_en), .Y(n1877)
         );
  INVX1 U2211 ( .A(n1878), .Y(n1359) );
  MUX2X1 U2212 ( .B(data_out[238]), .A(data_out[230]), .S(shift_en), .Y(n1878)
         );
  INVX1 U2213 ( .A(n1879), .Y(n1357) );
  MUX2X1 U2214 ( .B(data_out[246]), .A(data_out[238]), .S(shift_en), .Y(n1879)
         );
  INVX1 U2215 ( .A(n1880), .Y(n1355) );
  MUX2X1 U2216 ( .B(data_out[254]), .A(data_out[246]), .S(shift_en), .Y(n1880)
         );
  INVX1 U2217 ( .A(n1881), .Y(n1353) );
  MUX2X1 U2218 ( .B(data_out[262]), .A(data_out[254]), .S(shift_en), .Y(n1881)
         );
  INVX1 U2219 ( .A(n1882), .Y(n1351) );
  MUX2X1 U2220 ( .B(data_out[270]), .A(data_out[262]), .S(shift_en), .Y(n1882)
         );
  INVX1 U2221 ( .A(n1883), .Y(n1349) );
  MUX2X1 U2222 ( .B(data_out[278]), .A(data_out[270]), .S(shift_en), .Y(n1883)
         );
  INVX1 U2223 ( .A(n1884), .Y(n1347) );
  MUX2X1 U2224 ( .B(data_out[286]), .A(data_out[278]), .S(shift_en), .Y(n1884)
         );
  INVX1 U2225 ( .A(n1885), .Y(n1345) );
  MUX2X1 U2226 ( .B(data_out[294]), .A(data_out[286]), .S(shift_en), .Y(n1885)
         );
  INVX1 U2227 ( .A(n1886), .Y(n1343) );
  MUX2X1 U2228 ( .B(data_out[302]), .A(data_out[294]), .S(shift_en), .Y(n1886)
         );
  INVX1 U2229 ( .A(n1887), .Y(n1341) );
  MUX2X1 U2230 ( .B(data_out[310]), .A(data_out[302]), .S(shift_en), .Y(n1887)
         );
  INVX1 U2231 ( .A(n1888), .Y(n1339) );
  MUX2X1 U2232 ( .B(data_out[318]), .A(data_out[310]), .S(shift_en), .Y(n1888)
         );
  INVX1 U2233 ( .A(n1889), .Y(n1337) );
  MUX2X1 U2234 ( .B(data_out[326]), .A(data_out[318]), .S(shift_en), .Y(n1889)
         );
  INVX1 U2235 ( .A(n1890), .Y(n1335) );
  MUX2X1 U2236 ( .B(data_out[334]), .A(data_out[326]), .S(shift_en), .Y(n1890)
         );
  INVX1 U2237 ( .A(n1891), .Y(n1333) );
  MUX2X1 U2238 ( .B(data_out[342]), .A(data_out[334]), .S(shift_en), .Y(n1891)
         );
  INVX1 U2239 ( .A(n1892), .Y(n1331) );
  MUX2X1 U2240 ( .B(data_out[350]), .A(data_out[342]), .S(shift_en), .Y(n1892)
         );
  INVX1 U2241 ( .A(n1893), .Y(n1329) );
  MUX2X1 U2242 ( .B(data_out[358]), .A(data_out[350]), .S(shift_en), .Y(n1893)
         );
  INVX1 U2243 ( .A(n1894), .Y(n1327) );
  MUX2X1 U2244 ( .B(data_out[366]), .A(data_out[358]), .S(shift_en), .Y(n1894)
         );
  INVX1 U2245 ( .A(n1895), .Y(n1325) );
  MUX2X1 U2246 ( .B(data_out[374]), .A(data_out[366]), .S(shift_en), .Y(n1895)
         );
  INVX1 U2247 ( .A(n1896), .Y(n1323) );
  MUX2X1 U2248 ( .B(data_out[382]), .A(data_out[374]), .S(shift_en), .Y(n1896)
         );
  INVX1 U2249 ( .A(n1897), .Y(n1321) );
  MUX2X1 U2250 ( .B(data_out[390]), .A(data_out[382]), .S(shift_en), .Y(n1897)
         );
  INVX1 U2251 ( .A(n1898), .Y(n1319) );
  MUX2X1 U2252 ( .B(data_out[398]), .A(data_out[390]), .S(shift_en), .Y(n1898)
         );
  INVX1 U2253 ( .A(n1899), .Y(n1317) );
  MUX2X1 U2254 ( .B(data_out[406]), .A(data_out[398]), .S(shift_en), .Y(n1899)
         );
  INVX1 U2255 ( .A(n1900), .Y(n1315) );
  MUX2X1 U2256 ( .B(data_out[414]), .A(data_out[406]), .S(shift_en), .Y(n1900)
         );
  INVX1 U2257 ( .A(n1901), .Y(n1313) );
  MUX2X1 U2258 ( .B(data_out[422]), .A(data_out[414]), .S(shift_en), .Y(n1901)
         );
  INVX1 U2259 ( .A(n1902), .Y(n1311) );
  MUX2X1 U2260 ( .B(data_out[430]), .A(data_out[422]), .S(shift_en), .Y(n1902)
         );
  INVX1 U2261 ( .A(n1903), .Y(n1309) );
  MUX2X1 U2262 ( .B(data_out[438]), .A(data_out[430]), .S(shift_en), .Y(n1903)
         );
  INVX1 U2263 ( .A(n1904), .Y(n1307) );
  MUX2X1 U2264 ( .B(data_out[446]), .A(data_out[438]), .S(shift_en), .Y(n1904)
         );
  INVX1 U2265 ( .A(n1905), .Y(n1305) );
  MUX2X1 U2266 ( .B(data_out[454]), .A(data_out[446]), .S(shift_en), .Y(n1905)
         );
  INVX1 U2267 ( .A(n1906), .Y(n1303) );
  MUX2X1 U2268 ( .B(data_out[462]), .A(data_out[454]), .S(shift_en), .Y(n1906)
         );
  INVX1 U2269 ( .A(n1907), .Y(n1301) );
  MUX2X1 U2270 ( .B(data_out[470]), .A(data_out[462]), .S(shift_en), .Y(n1907)
         );
  INVX1 U2271 ( .A(n1908), .Y(n1299) );
  MUX2X1 U2272 ( .B(data_out[478]), .A(data_out[470]), .S(shift_en), .Y(n1908)
         );
  INVX1 U2273 ( .A(n1909), .Y(n1297) );
  MUX2X1 U2274 ( .B(data_out[486]), .A(data_out[478]), .S(shift_en), .Y(n1909)
         );
  INVX1 U2275 ( .A(n1910), .Y(n1295) );
  MUX2X1 U2276 ( .B(data_out[494]), .A(data_out[486]), .S(shift_en), .Y(n1910)
         );
  INVX1 U2277 ( .A(n1911), .Y(n1293) );
  MUX2X1 U2278 ( .B(data_out[502]), .A(data_out[494]), .S(shift_en), .Y(n1911)
         );
  INVX1 U2279 ( .A(n1912), .Y(n1291) );
  MUX2X1 U2280 ( .B(data_out[510]), .A(data_out[502]), .S(shift_en), .Y(n1912)
         );
  INVX1 U2281 ( .A(n1913), .Y(n1289) );
  MUX2X1 U2282 ( .B(data_out[5]), .A(data_in[5]), .S(shift_en), .Y(n1913) );
  INVX1 U2283 ( .A(n1914), .Y(n1287) );
  MUX2X1 U2284 ( .B(data_out[13]), .A(data_out[5]), .S(shift_en), .Y(n1914) );
  INVX1 U2285 ( .A(n1915), .Y(n1285) );
  MUX2X1 U2286 ( .B(data_out[21]), .A(data_out[13]), .S(shift_en), .Y(n1915)
         );
  INVX1 U2287 ( .A(n1916), .Y(n1283) );
  MUX2X1 U2288 ( .B(data_out[29]), .A(data_out[21]), .S(shift_en), .Y(n1916)
         );
  INVX1 U2289 ( .A(n1917), .Y(n1281) );
  MUX2X1 U2290 ( .B(data_out[37]), .A(data_out[29]), .S(shift_en), .Y(n1917)
         );
  INVX1 U2291 ( .A(n1918), .Y(n1279) );
  MUX2X1 U2292 ( .B(data_out[45]), .A(data_out[37]), .S(shift_en), .Y(n1918)
         );
  INVX1 U2293 ( .A(n1919), .Y(n1277) );
  MUX2X1 U2294 ( .B(data_out[53]), .A(data_out[45]), .S(shift_en), .Y(n1919)
         );
  INVX1 U2295 ( .A(n1920), .Y(n1275) );
  MUX2X1 U2296 ( .B(data_out[61]), .A(data_out[53]), .S(shift_en), .Y(n1920)
         );
  INVX1 U2297 ( .A(n1921), .Y(n1273) );
  MUX2X1 U2298 ( .B(data_out[69]), .A(data_out[61]), .S(shift_en), .Y(n1921)
         );
  INVX1 U2299 ( .A(n1922), .Y(n1271) );
  MUX2X1 U2300 ( .B(data_out[77]), .A(data_out[69]), .S(shift_en), .Y(n1922)
         );
  INVX1 U2301 ( .A(n1923), .Y(n1269) );
  MUX2X1 U2302 ( .B(data_out[85]), .A(data_out[77]), .S(shift_en), .Y(n1923)
         );
  INVX1 U2303 ( .A(n1924), .Y(n1267) );
  MUX2X1 U2304 ( .B(data_out[93]), .A(data_out[85]), .S(shift_en), .Y(n1924)
         );
  INVX1 U2305 ( .A(n1925), .Y(n1265) );
  MUX2X1 U2306 ( .B(data_out[101]), .A(data_out[93]), .S(shift_en), .Y(n1925)
         );
  INVX1 U2307 ( .A(n1926), .Y(n1263) );
  MUX2X1 U2308 ( .B(data_out[109]), .A(data_out[101]), .S(shift_en), .Y(n1926)
         );
  INVX1 U2309 ( .A(n1927), .Y(n1261) );
  MUX2X1 U2310 ( .B(data_out[117]), .A(data_out[109]), .S(shift_en), .Y(n1927)
         );
  INVX1 U2311 ( .A(n1928), .Y(n1259) );
  MUX2X1 U2312 ( .B(data_out[125]), .A(data_out[117]), .S(shift_en), .Y(n1928)
         );
  INVX1 U2313 ( .A(n1929), .Y(n1257) );
  MUX2X1 U2314 ( .B(data_out[133]), .A(data_out[125]), .S(shift_en), .Y(n1929)
         );
  INVX1 U2315 ( .A(n1930), .Y(n1255) );
  MUX2X1 U2316 ( .B(data_out[141]), .A(data_out[133]), .S(shift_en), .Y(n1930)
         );
  INVX1 U2317 ( .A(n1931), .Y(n1253) );
  MUX2X1 U2318 ( .B(data_out[149]), .A(data_out[141]), .S(shift_en), .Y(n1931)
         );
  INVX1 U2319 ( .A(n1932), .Y(n1251) );
  MUX2X1 U2320 ( .B(data_out[157]), .A(data_out[149]), .S(shift_en), .Y(n1932)
         );
  INVX1 U2321 ( .A(n1933), .Y(n1249) );
  MUX2X1 U2322 ( .B(data_out[165]), .A(data_out[157]), .S(shift_en), .Y(n1933)
         );
  INVX1 U2323 ( .A(n1934), .Y(n1247) );
  MUX2X1 U2324 ( .B(data_out[173]), .A(data_out[165]), .S(shift_en), .Y(n1934)
         );
  INVX1 U2325 ( .A(n1935), .Y(n1245) );
  MUX2X1 U2326 ( .B(data_out[181]), .A(data_out[173]), .S(shift_en), .Y(n1935)
         );
  INVX1 U2327 ( .A(n1936), .Y(n1243) );
  MUX2X1 U2328 ( .B(data_out[189]), .A(data_out[181]), .S(shift_en), .Y(n1936)
         );
  INVX1 U2329 ( .A(n1937), .Y(n1241) );
  MUX2X1 U2330 ( .B(data_out[197]), .A(data_out[189]), .S(shift_en), .Y(n1937)
         );
  INVX1 U2331 ( .A(n1938), .Y(n1239) );
  MUX2X1 U2332 ( .B(data_out[205]), .A(data_out[197]), .S(shift_en), .Y(n1938)
         );
  INVX1 U2333 ( .A(n1939), .Y(n1237) );
  MUX2X1 U2334 ( .B(data_out[213]), .A(data_out[205]), .S(shift_en), .Y(n1939)
         );
  INVX1 U2335 ( .A(n1940), .Y(n1235) );
  MUX2X1 U2336 ( .B(data_out[221]), .A(data_out[213]), .S(shift_en), .Y(n1940)
         );
  INVX1 U2337 ( .A(n1941), .Y(n1233) );
  MUX2X1 U2338 ( .B(data_out[229]), .A(data_out[221]), .S(shift_en), .Y(n1941)
         );
  INVX1 U2339 ( .A(n1942), .Y(n1231) );
  MUX2X1 U2340 ( .B(data_out[237]), .A(data_out[229]), .S(shift_en), .Y(n1942)
         );
  INVX1 U2341 ( .A(n1943), .Y(n1229) );
  MUX2X1 U2342 ( .B(data_out[245]), .A(data_out[237]), .S(shift_en), .Y(n1943)
         );
  INVX1 U2343 ( .A(n1944), .Y(n1227) );
  MUX2X1 U2344 ( .B(data_out[253]), .A(data_out[245]), .S(shift_en), .Y(n1944)
         );
  INVX1 U2345 ( .A(n1945), .Y(n1225) );
  MUX2X1 U2346 ( .B(data_out[261]), .A(data_out[253]), .S(shift_en), .Y(n1945)
         );
  INVX1 U2347 ( .A(n1946), .Y(n1223) );
  MUX2X1 U2348 ( .B(data_out[269]), .A(data_out[261]), .S(shift_en), .Y(n1946)
         );
  INVX1 U2349 ( .A(n1947), .Y(n1221) );
  MUX2X1 U2350 ( .B(data_out[277]), .A(data_out[269]), .S(shift_en), .Y(n1947)
         );
  INVX1 U2351 ( .A(n1948), .Y(n1219) );
  MUX2X1 U2352 ( .B(data_out[285]), .A(data_out[277]), .S(shift_en), .Y(n1948)
         );
  INVX1 U2353 ( .A(n1949), .Y(n1217) );
  MUX2X1 U2354 ( .B(data_out[293]), .A(data_out[285]), .S(shift_en), .Y(n1949)
         );
  INVX1 U2355 ( .A(n1950), .Y(n1215) );
  MUX2X1 U2356 ( .B(data_out[301]), .A(data_out[293]), .S(shift_en), .Y(n1950)
         );
  INVX1 U2357 ( .A(n1951), .Y(n1213) );
  MUX2X1 U2358 ( .B(data_out[309]), .A(data_out[301]), .S(shift_en), .Y(n1951)
         );
  INVX1 U2359 ( .A(n1952), .Y(n1211) );
  MUX2X1 U2360 ( .B(data_out[317]), .A(data_out[309]), .S(shift_en), .Y(n1952)
         );
  INVX1 U2361 ( .A(n1953), .Y(n1209) );
  MUX2X1 U2362 ( .B(data_out[325]), .A(data_out[317]), .S(shift_en), .Y(n1953)
         );
  INVX1 U2363 ( .A(n1954), .Y(n1207) );
  MUX2X1 U2364 ( .B(data_out[333]), .A(data_out[325]), .S(shift_en), .Y(n1954)
         );
  INVX1 U2365 ( .A(n1955), .Y(n1205) );
  MUX2X1 U2366 ( .B(data_out[341]), .A(data_out[333]), .S(shift_en), .Y(n1955)
         );
  INVX1 U2367 ( .A(n1956), .Y(n1203) );
  MUX2X1 U2368 ( .B(data_out[349]), .A(data_out[341]), .S(shift_en), .Y(n1956)
         );
  INVX1 U2369 ( .A(n1957), .Y(n1201) );
  MUX2X1 U2370 ( .B(data_out[357]), .A(data_out[349]), .S(shift_en), .Y(n1957)
         );
  INVX1 U2371 ( .A(n1958), .Y(n1199) );
  MUX2X1 U2372 ( .B(data_out[365]), .A(data_out[357]), .S(shift_en), .Y(n1958)
         );
  INVX1 U2373 ( .A(n1959), .Y(n1197) );
  MUX2X1 U2374 ( .B(data_out[373]), .A(data_out[365]), .S(shift_en), .Y(n1959)
         );
  INVX1 U2375 ( .A(n1960), .Y(n1195) );
  MUX2X1 U2376 ( .B(data_out[381]), .A(data_out[373]), .S(shift_en), .Y(n1960)
         );
  INVX1 U2377 ( .A(n1961), .Y(n1193) );
  MUX2X1 U2378 ( .B(data_out[389]), .A(data_out[381]), .S(shift_en), .Y(n1961)
         );
  INVX1 U2379 ( .A(n1962), .Y(n1191) );
  MUX2X1 U2380 ( .B(data_out[397]), .A(data_out[389]), .S(shift_en), .Y(n1962)
         );
  INVX1 U2381 ( .A(n1963), .Y(n1189) );
  MUX2X1 U2382 ( .B(data_out[405]), .A(data_out[397]), .S(shift_en), .Y(n1963)
         );
  INVX1 U2383 ( .A(n1964), .Y(n1187) );
  MUX2X1 U2384 ( .B(data_out[413]), .A(data_out[405]), .S(shift_en), .Y(n1964)
         );
  INVX1 U2385 ( .A(n1965), .Y(n1185) );
  MUX2X1 U2386 ( .B(data_out[421]), .A(data_out[413]), .S(shift_en), .Y(n1965)
         );
  INVX1 U2387 ( .A(n1966), .Y(n1183) );
  MUX2X1 U2388 ( .B(data_out[429]), .A(data_out[421]), .S(shift_en), .Y(n1966)
         );
  INVX1 U2389 ( .A(n1967), .Y(n1181) );
  MUX2X1 U2390 ( .B(data_out[437]), .A(data_out[429]), .S(shift_en), .Y(n1967)
         );
  INVX1 U2391 ( .A(n1968), .Y(n1179) );
  MUX2X1 U2392 ( .B(data_out[445]), .A(data_out[437]), .S(shift_en), .Y(n1968)
         );
  INVX1 U2393 ( .A(n1969), .Y(n1177) );
  MUX2X1 U2394 ( .B(data_out[453]), .A(data_out[445]), .S(shift_en), .Y(n1969)
         );
  INVX1 U2395 ( .A(n1970), .Y(n1175) );
  MUX2X1 U2396 ( .B(data_out[461]), .A(data_out[453]), .S(shift_en), .Y(n1970)
         );
  INVX1 U2397 ( .A(n1971), .Y(n1173) );
  MUX2X1 U2398 ( .B(data_out[469]), .A(data_out[461]), .S(shift_en), .Y(n1971)
         );
  INVX1 U2399 ( .A(n1972), .Y(n1171) );
  MUX2X1 U2400 ( .B(data_out[477]), .A(data_out[469]), .S(shift_en), .Y(n1972)
         );
  INVX1 U2401 ( .A(n1973), .Y(n1169) );
  MUX2X1 U2402 ( .B(data_out[485]), .A(data_out[477]), .S(shift_en), .Y(n1973)
         );
  INVX1 U2403 ( .A(n1974), .Y(n1167) );
  MUX2X1 U2404 ( .B(data_out[493]), .A(data_out[485]), .S(shift_en), .Y(n1974)
         );
  INVX1 U2405 ( .A(n1975), .Y(n1165) );
  MUX2X1 U2406 ( .B(data_out[501]), .A(data_out[493]), .S(shift_en), .Y(n1975)
         );
  INVX1 U2407 ( .A(n1976), .Y(n1163) );
  MUX2X1 U2408 ( .B(data_out[509]), .A(data_out[501]), .S(shift_en), .Y(n1976)
         );
  INVX1 U2409 ( .A(n1977), .Y(n1161) );
  MUX2X1 U2410 ( .B(data_out[4]), .A(data_in[4]), .S(shift_en), .Y(n1977) );
  INVX1 U2411 ( .A(n1978), .Y(n1159) );
  MUX2X1 U2412 ( .B(data_out[12]), .A(data_out[4]), .S(shift_en), .Y(n1978) );
  INVX1 U2413 ( .A(n1979), .Y(n1157) );
  MUX2X1 U2414 ( .B(data_out[20]), .A(data_out[12]), .S(shift_en), .Y(n1979)
         );
  INVX1 U2415 ( .A(n1980), .Y(n1155) );
  MUX2X1 U2416 ( .B(data_out[28]), .A(data_out[20]), .S(shift_en), .Y(n1980)
         );
  INVX1 U2417 ( .A(n1981), .Y(n1153) );
  MUX2X1 U2418 ( .B(data_out[36]), .A(data_out[28]), .S(shift_en), .Y(n1981)
         );
  INVX1 U2419 ( .A(n1982), .Y(n1151) );
  MUX2X1 U2420 ( .B(data_out[44]), .A(data_out[36]), .S(shift_en), .Y(n1982)
         );
  INVX1 U2421 ( .A(n1983), .Y(n1149) );
  MUX2X1 U2422 ( .B(data_out[52]), .A(data_out[44]), .S(shift_en), .Y(n1983)
         );
  INVX1 U2423 ( .A(n1984), .Y(n1147) );
  MUX2X1 U2424 ( .B(data_out[60]), .A(data_out[52]), .S(shift_en), .Y(n1984)
         );
  INVX1 U2425 ( .A(n1985), .Y(n1145) );
  MUX2X1 U2426 ( .B(data_out[68]), .A(data_out[60]), .S(shift_en), .Y(n1985)
         );
  INVX1 U2427 ( .A(n1986), .Y(n1143) );
  MUX2X1 U2428 ( .B(data_out[76]), .A(data_out[68]), .S(shift_en), .Y(n1986)
         );
  INVX1 U2429 ( .A(n1987), .Y(n1141) );
  MUX2X1 U2430 ( .B(data_out[84]), .A(data_out[76]), .S(shift_en), .Y(n1987)
         );
  INVX1 U2431 ( .A(n1988), .Y(n1139) );
  MUX2X1 U2432 ( .B(data_out[92]), .A(data_out[84]), .S(shift_en), .Y(n1988)
         );
  INVX1 U2433 ( .A(n1989), .Y(n1137) );
  MUX2X1 U2434 ( .B(data_out[100]), .A(data_out[92]), .S(shift_en), .Y(n1989)
         );
  INVX1 U2435 ( .A(n1990), .Y(n1135) );
  MUX2X1 U2436 ( .B(data_out[108]), .A(data_out[100]), .S(shift_en), .Y(n1990)
         );
  INVX1 U2437 ( .A(n1991), .Y(n1133) );
  MUX2X1 U2438 ( .B(data_out[116]), .A(data_out[108]), .S(shift_en), .Y(n1991)
         );
  INVX1 U2439 ( .A(n1992), .Y(n1131) );
  MUX2X1 U2440 ( .B(data_out[124]), .A(data_out[116]), .S(shift_en), .Y(n1992)
         );
  INVX1 U2441 ( .A(n1993), .Y(n1129) );
  MUX2X1 U2442 ( .B(data_out[132]), .A(data_out[124]), .S(shift_en), .Y(n1993)
         );
  INVX1 U2443 ( .A(n1994), .Y(n1127) );
  MUX2X1 U2444 ( .B(data_out[140]), .A(data_out[132]), .S(shift_en), .Y(n1994)
         );
  INVX1 U2445 ( .A(n1995), .Y(n1125) );
  MUX2X1 U2446 ( .B(data_out[148]), .A(data_out[140]), .S(shift_en), .Y(n1995)
         );
  INVX1 U2447 ( .A(n1996), .Y(n1123) );
  MUX2X1 U2448 ( .B(data_out[156]), .A(data_out[148]), .S(shift_en), .Y(n1996)
         );
  INVX1 U2449 ( .A(n1997), .Y(n1121) );
  MUX2X1 U2450 ( .B(data_out[164]), .A(data_out[156]), .S(shift_en), .Y(n1997)
         );
  INVX1 U2451 ( .A(n1998), .Y(n1119) );
  MUX2X1 U2452 ( .B(data_out[172]), .A(data_out[164]), .S(shift_en), .Y(n1998)
         );
  INVX1 U2453 ( .A(n1999), .Y(n1117) );
  MUX2X1 U2454 ( .B(data_out[180]), .A(data_out[172]), .S(shift_en), .Y(n1999)
         );
  INVX1 U2455 ( .A(n2000), .Y(n1115) );
  MUX2X1 U2456 ( .B(data_out[188]), .A(data_out[180]), .S(shift_en), .Y(n2000)
         );
  INVX1 U2457 ( .A(n2001), .Y(n1113) );
  MUX2X1 U2458 ( .B(data_out[196]), .A(data_out[188]), .S(shift_en), .Y(n2001)
         );
  INVX1 U2459 ( .A(n2002), .Y(n1111) );
  MUX2X1 U2460 ( .B(data_out[204]), .A(data_out[196]), .S(shift_en), .Y(n2002)
         );
  INVX1 U2461 ( .A(n2003), .Y(n1109) );
  MUX2X1 U2462 ( .B(data_out[212]), .A(data_out[204]), .S(shift_en), .Y(n2003)
         );
  INVX1 U2463 ( .A(n2004), .Y(n1107) );
  MUX2X1 U2464 ( .B(data_out[220]), .A(data_out[212]), .S(shift_en), .Y(n2004)
         );
  INVX1 U2465 ( .A(n2005), .Y(n1105) );
  MUX2X1 U2466 ( .B(data_out[228]), .A(data_out[220]), .S(shift_en), .Y(n2005)
         );
  INVX1 U2467 ( .A(n2006), .Y(n1103) );
  MUX2X1 U2468 ( .B(data_out[236]), .A(data_out[228]), .S(shift_en), .Y(n2006)
         );
  INVX1 U2469 ( .A(n2007), .Y(n1101) );
  MUX2X1 U2470 ( .B(data_out[244]), .A(data_out[236]), .S(shift_en), .Y(n2007)
         );
  INVX1 U2471 ( .A(n2008), .Y(n1099) );
  MUX2X1 U2472 ( .B(data_out[252]), .A(data_out[244]), .S(shift_en), .Y(n2008)
         );
  INVX1 U2473 ( .A(n2009), .Y(n1097) );
  MUX2X1 U2474 ( .B(data_out[260]), .A(data_out[252]), .S(shift_en), .Y(n2009)
         );
  INVX1 U2475 ( .A(n2010), .Y(n1095) );
  MUX2X1 U2476 ( .B(data_out[268]), .A(data_out[260]), .S(shift_en), .Y(n2010)
         );
  INVX1 U2477 ( .A(n2011), .Y(n1093) );
  MUX2X1 U2478 ( .B(data_out[276]), .A(data_out[268]), .S(shift_en), .Y(n2011)
         );
  INVX1 U2479 ( .A(n2012), .Y(n1091) );
  MUX2X1 U2480 ( .B(data_out[284]), .A(data_out[276]), .S(shift_en), .Y(n2012)
         );
  INVX1 U2481 ( .A(n2013), .Y(n1089) );
  MUX2X1 U2482 ( .B(data_out[292]), .A(data_out[284]), .S(shift_en), .Y(n2013)
         );
  INVX1 U2483 ( .A(n2014), .Y(n1087) );
  MUX2X1 U2484 ( .B(data_out[300]), .A(data_out[292]), .S(shift_en), .Y(n2014)
         );
  INVX1 U2485 ( .A(n2015), .Y(n1085) );
  MUX2X1 U2486 ( .B(data_out[308]), .A(data_out[300]), .S(shift_en), .Y(n2015)
         );
  INVX1 U2487 ( .A(n2016), .Y(n1083) );
  MUX2X1 U2488 ( .B(data_out[316]), .A(data_out[308]), .S(shift_en), .Y(n2016)
         );
  INVX1 U2489 ( .A(n2017), .Y(n1081) );
  MUX2X1 U2490 ( .B(data_out[324]), .A(data_out[316]), .S(shift_en), .Y(n2017)
         );
  INVX1 U2491 ( .A(n2018), .Y(n1079) );
  MUX2X1 U2492 ( .B(data_out[332]), .A(data_out[324]), .S(shift_en), .Y(n2018)
         );
  INVX1 U2493 ( .A(n2019), .Y(n1077) );
  MUX2X1 U2494 ( .B(data_out[340]), .A(data_out[332]), .S(shift_en), .Y(n2019)
         );
  INVX1 U2495 ( .A(n2020), .Y(n1075) );
  MUX2X1 U2496 ( .B(data_out[348]), .A(data_out[340]), .S(shift_en), .Y(n2020)
         );
  INVX1 U2497 ( .A(n2021), .Y(n1073) );
  MUX2X1 U2498 ( .B(data_out[356]), .A(data_out[348]), .S(shift_en), .Y(n2021)
         );
  INVX1 U2499 ( .A(n2022), .Y(n1071) );
  MUX2X1 U2500 ( .B(data_out[364]), .A(data_out[356]), .S(shift_en), .Y(n2022)
         );
  INVX1 U2501 ( .A(n2023), .Y(n1069) );
  MUX2X1 U2502 ( .B(data_out[372]), .A(data_out[364]), .S(shift_en), .Y(n2023)
         );
  INVX1 U2503 ( .A(n2024), .Y(n1067) );
  MUX2X1 U2504 ( .B(data_out[380]), .A(data_out[372]), .S(shift_en), .Y(n2024)
         );
  INVX1 U2505 ( .A(n2025), .Y(n1065) );
  MUX2X1 U2506 ( .B(data_out[388]), .A(data_out[380]), .S(shift_en), .Y(n2025)
         );
  INVX1 U2507 ( .A(n2026), .Y(n1063) );
  MUX2X1 U2508 ( .B(data_out[396]), .A(data_out[388]), .S(shift_en), .Y(n2026)
         );
  INVX1 U2509 ( .A(n2027), .Y(n1061) );
  MUX2X1 U2510 ( .B(data_out[404]), .A(data_out[396]), .S(shift_en), .Y(n2027)
         );
  INVX1 U2511 ( .A(n2028), .Y(n1059) );
  MUX2X1 U2512 ( .B(data_out[412]), .A(data_out[404]), .S(shift_en), .Y(n2028)
         );
  INVX1 U2513 ( .A(n2029), .Y(n1057) );
  MUX2X1 U2514 ( .B(data_out[420]), .A(data_out[412]), .S(shift_en), .Y(n2029)
         );
  INVX1 U2515 ( .A(n2030), .Y(n1055) );
  MUX2X1 U2516 ( .B(data_out[428]), .A(data_out[420]), .S(shift_en), .Y(n2030)
         );
  INVX1 U2517 ( .A(n2031), .Y(n1053) );
  MUX2X1 U2518 ( .B(data_out[436]), .A(data_out[428]), .S(shift_en), .Y(n2031)
         );
  INVX1 U2519 ( .A(n2032), .Y(n1051) );
  MUX2X1 U2520 ( .B(data_out[444]), .A(data_out[436]), .S(shift_en), .Y(n2032)
         );
  INVX1 U2521 ( .A(n2033), .Y(n1049) );
  MUX2X1 U2522 ( .B(data_out[452]), .A(data_out[444]), .S(shift_en), .Y(n2033)
         );
  INVX1 U2523 ( .A(n2034), .Y(n1047) );
  MUX2X1 U2524 ( .B(data_out[460]), .A(data_out[452]), .S(shift_en), .Y(n2034)
         );
  INVX1 U2525 ( .A(n2035), .Y(n1045) );
  MUX2X1 U2526 ( .B(data_out[468]), .A(data_out[460]), .S(shift_en), .Y(n2035)
         );
  INVX1 U2527 ( .A(n2036), .Y(n1043) );
  MUX2X1 U2528 ( .B(data_out[476]), .A(data_out[468]), .S(shift_en), .Y(n2036)
         );
  INVX1 U2529 ( .A(n2037), .Y(n1041) );
  MUX2X1 U2530 ( .B(data_out[484]), .A(data_out[476]), .S(shift_en), .Y(n2037)
         );
  INVX1 U2531 ( .A(n2038), .Y(n1039) );
  MUX2X1 U2532 ( .B(data_out[492]), .A(data_out[484]), .S(shift_en), .Y(n2038)
         );
  INVX1 U2533 ( .A(n2039), .Y(n1037) );
  MUX2X1 U2534 ( .B(data_out[500]), .A(data_out[492]), .S(shift_en), .Y(n2039)
         );
  INVX1 U2535 ( .A(n2040), .Y(n1035) );
  MUX2X1 U2536 ( .B(data_out[508]), .A(data_out[500]), .S(shift_en), .Y(n2040)
         );
  INVX1 U2537 ( .A(n2041), .Y(n1033) );
  MUX2X1 U2538 ( .B(data_out[3]), .A(data_in[3]), .S(shift_en), .Y(n2041) );
  INVX1 U2539 ( .A(n2042), .Y(n1031) );
  MUX2X1 U2540 ( .B(data_out[11]), .A(data_out[3]), .S(shift_en), .Y(n2042) );
  INVX1 U2541 ( .A(n2043), .Y(n1029) );
  MUX2X1 U2542 ( .B(data_out[19]), .A(data_out[11]), .S(shift_en), .Y(n2043)
         );
  INVX1 U2543 ( .A(n2044), .Y(n1027) );
  MUX2X1 U2544 ( .B(data_out[27]), .A(data_out[19]), .S(shift_en), .Y(n2044)
         );
  INVX1 U2545 ( .A(n2045), .Y(n1025) );
  MUX2X1 U2546 ( .B(data_out[35]), .A(data_out[27]), .S(shift_en), .Y(n2045)
         );
  INVX1 U2547 ( .A(n2046), .Y(n1023) );
  MUX2X1 U2548 ( .B(data_out[43]), .A(data_out[35]), .S(shift_en), .Y(n2046)
         );
  INVX1 U2549 ( .A(n2047), .Y(n1021) );
  MUX2X1 U2550 ( .B(data_out[51]), .A(data_out[43]), .S(shift_en), .Y(n2047)
         );
  INVX1 U2551 ( .A(n2048), .Y(n1019) );
  MUX2X1 U2552 ( .B(data_out[59]), .A(data_out[51]), .S(shift_en), .Y(n2048)
         );
  INVX1 U2553 ( .A(n2049), .Y(n1017) );
  MUX2X1 U2554 ( .B(data_out[67]), .A(data_out[59]), .S(shift_en), .Y(n2049)
         );
  INVX1 U2555 ( .A(n2050), .Y(n1015) );
  MUX2X1 U2556 ( .B(data_out[75]), .A(data_out[67]), .S(shift_en), .Y(n2050)
         );
  INVX1 U2557 ( .A(n2051), .Y(n1013) );
  MUX2X1 U2558 ( .B(data_out[83]), .A(data_out[75]), .S(shift_en), .Y(n2051)
         );
  INVX1 U2559 ( .A(n2052), .Y(n1011) );
  MUX2X1 U2560 ( .B(data_out[91]), .A(data_out[83]), .S(shift_en), .Y(n2052)
         );
  INVX1 U2561 ( .A(n2053), .Y(n1009) );
  MUX2X1 U2562 ( .B(data_out[99]), .A(data_out[91]), .S(shift_en), .Y(n2053)
         );
  INVX1 U2563 ( .A(n2054), .Y(n1007) );
  MUX2X1 U2564 ( .B(data_out[107]), .A(data_out[99]), .S(shift_en), .Y(n2054)
         );
  INVX1 U2565 ( .A(n2055), .Y(n1005) );
  MUX2X1 U2566 ( .B(data_out[115]), .A(data_out[107]), .S(shift_en), .Y(n2055)
         );
  INVX1 U2567 ( .A(n2056), .Y(n1003) );
  MUX2X1 U2568 ( .B(data_out[123]), .A(data_out[115]), .S(shift_en), .Y(n2056)
         );
  INVX1 U2569 ( .A(n2057), .Y(n1001) );
  MUX2X1 U2570 ( .B(data_out[131]), .A(data_out[123]), .S(shift_en), .Y(n2057)
         );
endmodule

