// $Id: $
// File name:   tb_usb_crc16.sv
// Created:     4/21/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: CRC16 testbench

`timescale 1ns / 10ps

module tb_usb_crc16_valid();
	
endmodule