// $Id: $
// File name:   datapath.sv
// Created:     4/16/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: Module for datapath block (interfaces with SRAM.
// 

module datapath
	(
		input [6:0] address_one,
		input [6:0] address_two,
		input [31:0] data_in,
		input [1:0] op_code,
		output [31:0] data_out
	);

endmodule