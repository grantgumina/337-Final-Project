// $Id: $
// File name:   usb_state_machine.sv
// Created:     4/16/2014
// Author:      Grant Gumina
// Lab Section: 02
// Version:     1.0  Initial Design Entry
// Description: USB Protocol State Machine

module usb_state_machine
	(
		input wire shift_out,
		input wire [7,0] data_in,
		output wire new_byte,
		output wire [7:0] data_out

		// OUTPUT WIRE USB DATA BUS??????
	);

endmodule